/////////////////////////////////////////////////////////////////////
////  AHB DMA Priority Encoder Sub-Module                        ////
////                                                             ////
////  Author: Ibrahim Hossam                                     ////
/////////////////////////////////////////////////////////////////////
module ahb_dma_pri_enc_sub(
valid,
pri_in,
pri_out);
//==========================================================================
// Inputs & Outputs
//==========================================================================
input		    valid;
input	[2:0]	pri_in;
output	[7:0]	pri_out;
//==========================================================================
// Internal signls
//==========================================================================
	reg	[7:0]	pri_out;
//==========================================================================
// Main code
//==========================================================================
	always_comb
	begin
		pri_out = (8'b1 << ({3{valid}} & pri_in));
	end

endmodule

