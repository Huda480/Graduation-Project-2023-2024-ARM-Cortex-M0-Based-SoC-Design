/////////////////////////////////////////////////////////////////////
////  AHB DMA oring array                                        ////
////                                                             ////
////  Author: Ibrahim Hossam                                     ////
/////////////////////////////////////////////////////////////////////
module or_opt #(
//==========================================================================
// Parameters
//==========================================================================
parameter channel_number = 15,width=5)(
//==========================================================================
// Inputs & Outputs
//==========================================================================
input   [width-1:0]     signals [0:channel_number-1] ,
output  [width-1:0]     ored_signal
);
//==========================================================================
// Internal signals
//==========================================================================
  reg     [width-1:0] ored_r  ;
//==========================================================================
// Main code
//==========================================================================
  always_comb begin
    ored_r = 8'h00; 
    foreach (signals[i]) begin
      ored_r |= signals[i]; 
    end
  end

  assign  ored_signal = ored_r;

endmodule