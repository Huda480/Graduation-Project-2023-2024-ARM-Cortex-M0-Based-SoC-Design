//==============================================================================
// Purpose: UART APB peripheral header
// Used in: cmsdk_apb_uart
//==============================================================================

// UART reset macros
`define ARM_UARTCTRL_RESET          10'b000
`define ARM_UARTBAUDDIV_RESET       20'b000