//==============================================================================
// Purpose: AHB slaves package
// Used in: cmsdk_iop_gpio
//==============================================================================
package ahb_pkg;
  //============================================================================
    //Include new data types
  //============================================================================
  typedef enum bit [1:0] 
  {
    IDLE      = 2'b00, 
    NOT_READY = 2'b10, 
    ERROR     = 2'b11
  } states_t;
  //============================================================================
endpackage: ahb_pkg