package compression_package;
localparam logic signed [1:0] Phi_var [96][64] = '{
		'{ 2'b01, 2'b00, 2'b00, 2'b01, 2'b01, 2'b01, 2'b11, 2'b00, 2'b10, 2'b00, 2'b01, 2'b00, 2'b00, 2'b00, 2'b11, 2'b00, 2'b01, 2'b10, 2'b11, 2'b00, 2'b00, 2'b00, 2'b01, 2'b01, 2'b00, 2'b11, 2'b00, 2'b11, 2'b11, 2'b00, 2'b10, 2'b01, 2'b01, 2'b10, 2'b00, 2'b11, 2'b00, 2'b00, 2'b01, 2'b00, 2'b01, 2'b00, 2'b00, 2'b01, 2'b01, 2'b01, 2'b11, 2'b11, 2'b01, 2'b00, 2'b10, 2'b10, 2'b00, 2'b00, 2'b00, 2'b11, 2'b01, 2'b01, 2'b00, 2'b01, 2'b11, 2'b00, 2'b10, 2'b11 },
		'{ 2'b11, 2'b00, 2'b01, 2'b10, 2'b00, 2'b01, 2'b00, 2'b11, 2'b00, 2'b01, 2'b10, 2'b01, 2'b11, 2'b00, 2'b00, 2'b00, 2'b01, 2'b11, 2'b10, 2'b00, 2'b00, 2'b11, 2'b00, 2'b00, 2'b10, 2'b11, 2'b00, 2'b00, 2'b10, 2'b11, 2'b00, 2'b00, 2'b01, 2'b11, 2'b10, 2'b11, 2'b00, 2'b00, 2'b00, 2'b11, 2'b01, 2'b00, 2'b01, 2'b01, 2'b11, 2'b10, 2'b11, 2'b00, 2'b00, 2'b01, 2'b10, 2'b01, 2'b01, 2'b01, 2'b11, 2'b11, 2'b01, 2'b01, 2'b00, 2'b01, 2'b11, 2'b00, 2'b11, 2'b00 },
		'{ 2'b01, 2'b11, 2'b11, 2'b00, 2'b01, 2'b11, 2'b00, 2'b00, 2'b00, 2'b01, 2'b00, 2'b00, 2'b11, 2'b01, 2'b00, 2'b00, 2'b10, 2'b00, 2'b01, 2'b11, 2'b10, 2'b11, 2'b10, 2'b00, 2'b00, 2'b01, 2'b11, 2'b01, 2'b00, 2'b00, 2'b11, 2'b00, 2'b11, 2'b00, 2'b00, 2'b00, 2'b11, 2'b10, 2'b11, 2'b00, 2'b00, 2'b00, 2'b10, 2'b01, 2'b00, 2'b01, 2'b00, 2'b11, 2'b01, 2'b00, 2'b00, 2'b00, 2'b00, 2'b11, 2'b11, 2'b01, 2'b10, 2'b01, 2'b01, 2'b11, 2'b00, 2'b11, 2'b11, 2'b11 },
		'{ 2'b00, 2'b11, 2'b00, 2'b01, 2'b11, 2'b00, 2'b00, 2'b01, 2'b11, 2'b01, 2'b00, 2'b11, 2'b00, 2'b11, 2'b11, 2'b01, 2'b01, 2'b00, 2'b01, 2'b00, 2'b00, 2'b01, 2'b01, 2'b00, 2'b00, 2'b00, 2'b01, 2'b00, 2'b11, 2'b00, 2'b00, 2'b00, 2'b11, 2'b10, 2'b00, 2'b00, 2'b11, 2'b00, 2'b11, 2'b10, 2'b01, 2'b00, 2'b00, 2'b11, 2'b00, 2'b01, 2'b00, 2'b01, 2'b11, 2'b01, 2'b00, 2'b01, 2'b10, 2'b01, 2'b10, 2'b00, 2'b01, 2'b01, 2'b10, 2'b01, 2'b11, 2'b01, 2'b11, 2'b00 },
		'{ 2'b00, 2'b11, 2'b01, 2'b11, 2'b01, 2'b11, 2'b00, 2'b01, 2'b00, 2'b01, 2'b00, 2'b01, 2'b00, 2'b01, 2'b01, 2'b11, 2'b01, 2'b00, 2'b01, 2'b01, 2'b10, 2'b10, 2'b01, 2'b00, 2'b00, 2'b00, 2'b00, 2'b01, 2'b11, 2'b00, 2'b01, 2'b00, 2'b11, 2'b11, 2'b01, 2'b00, 2'b00, 2'b00, 2'b11, 2'b01, 2'b01, 2'b01, 2'b11, 2'b11, 2'b01, 2'b11, 2'b00, 2'b00, 2'b01, 2'b11, 2'b11, 2'b01, 2'b00, 2'b11, 2'b01, 2'b11, 2'b01, 2'b00, 2'b10, 2'b01, 2'b01, 2'b11, 2'b00, 2'b01 },
		'{ 2'b00, 2'b11, 2'b10, 2'b00, 2'b10, 2'b11, 2'b00, 2'b00, 2'b00, 2'b10, 2'b11, 2'b01, 2'b00, 2'b01, 2'b01, 2'b10, 2'b00, 2'b01, 2'b00, 2'b11, 2'b01, 2'b00, 2'b00, 2'b00, 2'b00, 2'b01, 2'b01, 2'b11, 2'b11, 2'b01, 2'b01, 2'b11, 2'b11, 2'b00, 2'b01, 2'b00, 2'b01, 2'b01, 2'b01, 2'b00, 2'b11, 2'b00, 2'b00, 2'b11, 2'b01, 2'b00, 2'b00, 2'b11, 2'b11, 2'b11, 2'b00, 2'b00, 2'b01, 2'b00, 2'b01, 2'b01, 2'b00, 2'b11, 2'b01, 2'b00, 2'b11, 2'b11, 2'b11, 2'b01 },
		'{ 2'b01, 2'b00, 2'b01, 2'b00, 2'b01, 2'b01, 2'b10, 2'b01, 2'b00, 2'b00, 2'b00, 2'b10, 2'b11, 2'b00, 2'b00, 2'b11, 2'b00, 2'b01, 2'b01, 2'b10, 2'b00, 2'b00, 2'b11, 2'b11, 2'b00, 2'b00, 2'b01, 2'b00, 2'b10, 2'b01, 2'b01, 2'b11, 2'b01, 2'b01, 2'b11, 2'b01, 2'b11, 2'b11, 2'b00, 2'b01, 2'b00, 2'b11, 2'b00, 2'b00, 2'b00, 2'b11, 2'b00, 2'b11, 2'b00, 2'b01, 2'b00, 2'b00, 2'b10, 2'b01, 2'b00, 2'b00, 2'b00, 2'b00, 2'b01, 2'b00, 2'b10, 2'b01, 2'b01, 2'b11 },
		'{ 2'b01, 2'b11, 2'b01, 2'b11, 2'b00, 2'b11, 2'b11, 2'b00, 2'b00, 2'b00, 2'b01, 2'b11, 2'b00, 2'b01, 2'b01, 2'b11, 2'b00, 2'b11, 2'b01, 2'b01, 2'b00, 2'b01, 2'b01, 2'b11, 2'b01, 2'b01, 2'b00, 2'b10, 2'b00, 2'b01, 2'b01, 2'b00, 2'b11, 2'b00, 2'b01, 2'b01, 2'b00, 2'b01, 2'b00, 2'b11, 2'b11, 2'b11, 2'b11, 2'b00, 2'b01, 2'b00, 2'b10, 2'b00, 2'b01, 2'b00, 2'b01, 2'b10, 2'b00, 2'b01, 2'b00, 2'b00, 2'b11, 2'b01, 2'b10, 2'b11, 2'b00, 2'b01, 2'b01, 2'b11 },
		'{ 2'b01, 2'b11, 2'b01, 2'b11, 2'b00, 2'b01, 2'b11, 2'b10, 2'b00, 2'b00, 2'b01, 2'b11, 2'b01, 2'b01, 2'b11, 2'b00, 2'b10, 2'b01, 2'b01, 2'b00, 2'b11, 2'b10, 2'b01, 2'b00, 2'b01, 2'b01, 2'b00, 2'b00, 2'b01, 2'b00, 2'b00, 2'b00, 2'b01, 2'b11, 2'b11, 2'b01, 2'b11, 2'b11, 2'b00, 2'b10, 2'b11, 2'b00, 2'b11, 2'b01, 2'b00, 2'b00, 2'b01, 2'b10, 2'b00, 2'b00, 2'b00, 2'b11, 2'b01, 2'b00, 2'b00, 2'b11, 2'b00, 2'b01, 2'b01, 2'b01, 2'b00, 2'b01, 2'b01, 2'b10 },
		'{ 2'b11, 2'b01, 2'b00, 2'b00, 2'b00, 2'b10, 2'b11, 2'b00, 2'b00, 2'b11, 2'b01, 2'b10, 2'b00, 2'b00, 2'b10, 2'b01, 2'b00, 2'b11, 2'b01, 2'b00, 2'b11, 2'b00, 2'b11, 2'b01, 2'b01, 2'b11, 2'b01, 2'b11, 2'b00, 2'b11, 2'b00, 2'b11, 2'b00, 2'b11, 2'b00, 2'b11, 2'b00, 2'b11, 2'b11, 2'b00, 2'b00, 2'b01, 2'b11, 2'b01, 2'b11, 2'b01, 2'b00, 2'b00, 2'b00, 2'b00, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b11, 2'b00, 2'b11, 2'b10, 2'b00, 2'b11, 2'b11, 2'b01, 2'b11 },
		'{ 2'b01, 2'b00, 2'b01, 2'b00, 2'b00, 2'b00, 2'b01, 2'b01, 2'b01, 2'b11, 2'b00, 2'b01, 2'b11, 2'b00, 2'b00, 2'b00, 2'b00, 2'b00, 2'b01, 2'b11, 2'b00, 2'b00, 2'b00, 2'b11, 2'b00, 2'b01, 2'b01, 2'b01, 2'b01, 2'b00, 2'b11, 2'b00, 2'b11, 2'b01, 2'b00, 2'b00, 2'b10, 2'b01, 2'b11, 2'b00, 2'b01, 2'b01, 2'b00, 2'b10, 2'b01, 2'b01, 2'b01, 2'b11, 2'b00, 2'b11, 2'b01, 2'b01, 2'b01, 2'b11, 2'b00, 2'b00, 2'b11, 2'b00, 2'b10, 2'b00, 2'b01, 2'b00, 2'b00, 2'b11 },
		'{ 2'b11, 2'b00, 2'b01, 2'b01, 2'b00, 2'b00, 2'b01, 2'b00, 2'b01, 2'b01, 2'b10, 2'b10, 2'b00, 2'b00, 2'b00, 2'b00, 2'b00, 2'b11, 2'b00, 2'b00, 2'b00, 2'b01, 2'b01, 2'b10, 2'b00, 2'b01, 2'b01, 2'b01, 2'b00, 2'b11, 2'b00, 2'b00, 2'b10, 2'b00, 2'b01, 2'b11, 2'b00, 2'b00, 2'b11, 2'b01, 2'b11, 2'b11, 2'b00, 2'b10, 2'b10, 2'b11, 2'b00, 2'b01, 2'b11, 2'b00, 2'b01, 2'b11, 2'b11, 2'b10, 2'b01, 2'b11, 2'b01, 2'b01, 2'b00, 2'b00, 2'b11, 2'b01, 2'b00, 2'b00 },
		'{ 2'b11, 2'b00, 2'b11, 2'b01, 2'b01, 2'b01, 2'b11, 2'b00, 2'b00, 2'b00, 2'b11, 2'b11, 2'b11, 2'b11, 2'b00, 2'b11, 2'b00, 2'b11, 2'b01, 2'b00, 2'b10, 2'b00, 2'b00, 2'b11, 2'b00, 2'b00, 2'b01, 2'b00, 2'b00, 2'b11, 2'b10, 2'b11, 2'b00, 2'b01, 2'b11, 2'b00, 2'b00, 2'b01, 2'b00, 2'b00, 2'b01, 2'b11, 2'b00, 2'b01, 2'b11, 2'b11, 2'b11, 2'b00, 2'b10, 2'b00, 2'b01, 2'b01, 2'b01, 2'b11, 2'b11, 2'b10, 2'b01, 2'b01, 2'b11, 2'b00, 2'b00, 2'b11, 2'b01, 2'b01 },
		'{ 2'b01, 2'b11, 2'b00, 2'b11, 2'b01, 2'b01, 2'b11, 2'b01, 2'b01, 2'b11, 2'b11, 2'b00, 2'b11, 2'b00, 2'b00, 2'b00, 2'b00, 2'b00, 2'b00, 2'b11, 2'b00, 2'b01, 2'b00, 2'b01, 2'b00, 2'b00, 2'b11, 2'b11, 2'b00, 2'b01, 2'b10, 2'b00, 2'b11, 2'b01, 2'b11, 2'b10, 2'b00, 2'b00, 2'b10, 2'b01, 2'b01, 2'b11, 2'b01, 2'b00, 2'b00, 2'b01, 2'b11, 2'b11, 2'b00, 2'b00, 2'b00, 2'b10, 2'b01, 2'b01, 2'b00, 2'b00, 2'b00, 2'b01, 2'b11, 2'b01, 2'b00, 2'b01, 2'b01, 2'b11 },
		'{ 2'b01, 2'b00, 2'b10, 2'b01, 2'b00, 2'b01, 2'b01, 2'b11, 2'b00, 2'b00, 2'b01, 2'b00, 2'b01, 2'b00, 2'b01, 2'b00, 2'b01, 2'b11, 2'b01, 2'b11, 2'b00, 2'b11, 2'b00, 2'b01, 2'b01, 2'b01, 2'b01, 2'b10, 2'b00, 2'b00, 2'b01, 2'b01, 2'b00, 2'b00, 2'b00, 2'b00, 2'b00, 2'b01, 2'b11, 2'b01, 2'b00, 2'b11, 2'b11, 2'b00, 2'b00, 2'b10, 2'b01, 2'b00, 2'b01, 2'b01, 2'b01, 2'b01, 2'b10, 2'b00, 2'b00, 2'b11, 2'b11, 2'b00, 2'b10, 2'b00, 2'b01, 2'b11, 2'b00, 2'b00 },
		'{ 2'b01, 2'b01, 2'b01, 2'b00, 2'b00, 2'b01, 2'b00, 2'b11, 2'b00, 2'b01, 2'b11, 2'b01, 2'b01, 2'b11, 2'b00, 2'b11, 2'b11, 2'b11, 2'b00, 2'b01, 2'b11, 2'b11, 2'b00, 2'b11, 2'b01, 2'b01, 2'b11, 2'b00, 2'b11, 2'b00, 2'b01, 2'b01, 2'b10, 2'b00, 2'b01, 2'b00, 2'b11, 2'b00, 2'b01, 2'b01, 2'b00, 2'b00, 2'b11, 2'b11, 2'b00, 2'b00, 2'b11, 2'b11, 2'b01, 2'b00, 2'b01, 2'b01, 2'b01, 2'b01, 2'b00, 2'b01, 2'b00, 2'b01, 2'b11, 2'b00, 2'b11, 2'b10, 2'b10, 2'b01 },
		'{ 2'b11, 2'b01, 2'b00, 2'b00, 2'b11, 2'b00, 2'b00, 2'b01, 2'b01, 2'b01, 2'b11, 2'b00, 2'b00, 2'b01, 2'b00, 2'b00, 2'b11, 2'b11, 2'b01, 2'b01, 2'b01, 2'b00, 2'b11, 2'b01, 2'b11, 2'b01, 2'b11, 2'b00, 2'b01, 2'b01, 2'b01, 2'b01, 2'b11, 2'b11, 2'b01, 2'b00, 2'b01, 2'b01, 2'b00, 2'b01, 2'b10, 2'b00, 2'b11, 2'b11, 2'b10, 2'b11, 2'b01, 2'b11, 2'b01, 2'b00, 2'b00, 2'b01, 2'b01, 2'b01, 2'b10, 2'b00, 2'b01, 2'b00, 2'b11, 2'b11, 2'b11, 2'b10, 2'b11, 2'b01 },
		'{ 2'b11, 2'b01, 2'b11, 2'b10, 2'b11, 2'b00, 2'b01, 2'b00, 2'b01, 2'b00, 2'b00, 2'b01, 2'b00, 2'b11, 2'b01, 2'b01, 2'b11, 2'b00, 2'b01, 2'b00, 2'b00, 2'b00, 2'b01, 2'b00, 2'b01, 2'b01, 2'b01, 2'b00, 2'b01, 2'b11, 2'b11, 2'b11, 2'b00, 2'b01, 2'b00, 2'b10, 2'b00, 2'b00, 2'b11, 2'b11, 2'b10, 2'b01, 2'b00, 2'b01, 2'b01, 2'b01, 2'b11, 2'b01, 2'b00, 2'b00, 2'b01, 2'b00, 2'b01, 2'b01, 2'b10, 2'b11, 2'b01, 2'b00, 2'b00, 2'b10, 2'b11, 2'b01, 2'b11, 2'b11 },
		'{ 2'b11, 2'b01, 2'b01, 2'b00, 2'b11, 2'b01, 2'b01, 2'b01, 2'b01, 2'b11, 2'b11, 2'b01, 2'b00, 2'b00, 2'b11, 2'b01, 2'b01, 2'b00, 2'b00, 2'b01, 2'b11, 2'b00, 2'b01, 2'b00, 2'b00, 2'b01, 2'b11, 2'b00, 2'b11, 2'b10, 2'b11, 2'b11, 2'b00, 2'b00, 2'b01, 2'b00, 2'b01, 2'b10, 2'b11, 2'b00, 2'b11, 2'b01, 2'b10, 2'b01, 2'b10, 2'b01, 2'b00, 2'b01, 2'b01, 2'b11, 2'b00, 2'b11, 2'b00, 2'b10, 2'b01, 2'b00, 2'b00, 2'b00, 2'b00, 2'b10, 2'b01, 2'b10, 2'b10, 2'b01 },
		'{ 2'b11, 2'b00, 2'b10, 2'b00, 2'b00, 2'b01, 2'b00, 2'b11, 2'b00, 2'b11, 2'b00, 2'b10, 2'b01, 2'b00, 2'b00, 2'b00, 2'b11, 2'b00, 2'b00, 2'b01, 2'b00, 2'b11, 2'b00, 2'b01, 2'b01, 2'b00, 2'b11, 2'b00, 2'b01, 2'b01, 2'b00, 2'b11, 2'b01, 2'b00, 2'b11, 2'b11, 2'b01, 2'b00, 2'b01, 2'b01, 2'b00, 2'b11, 2'b00, 2'b11, 2'b11, 2'b00, 2'b01, 2'b11, 2'b11, 2'b00, 2'b01, 2'b11, 2'b01, 2'b10, 2'b01, 2'b01, 2'b01, 2'b00, 2'b01, 2'b00, 2'b00, 2'b11, 2'b01, 2'b00 },
		'{ 2'b11, 2'b11, 2'b00, 2'b00, 2'b00, 2'b10, 2'b10, 2'b11, 2'b00, 2'b01, 2'b01, 2'b01, 2'b01, 2'b11, 2'b00, 2'b01, 2'b01, 2'b00, 2'b00, 2'b00, 2'b11, 2'b10, 2'b01, 2'b00, 2'b00, 2'b10, 2'b11, 2'b01, 2'b01, 2'b11, 2'b11, 2'b01, 2'b00, 2'b11, 2'b00, 2'b00, 2'b01, 2'b01, 2'b01, 2'b00, 2'b10, 2'b01, 2'b11, 2'b11, 2'b01, 2'b00, 2'b00, 2'b01, 2'b11, 2'b01, 2'b00, 2'b00, 2'b00, 2'b01, 2'b00, 2'b11, 2'b00, 2'b00, 2'b00, 2'b11, 2'b11, 2'b01, 2'b00, 2'b00 },
		'{ 2'b11, 2'b10, 2'b01, 2'b00, 2'b11, 2'b00, 2'b10, 2'b11, 2'b11, 2'b10, 2'b11, 2'b00, 2'b00, 2'b01, 2'b00, 2'b01, 2'b00, 2'b00, 2'b00, 2'b01, 2'b00, 2'b01, 2'b01, 2'b11, 2'b00, 2'b01, 2'b00, 2'b00, 2'b11, 2'b01, 2'b01, 2'b00, 2'b00, 2'b00, 2'b10, 2'b10, 2'b10, 2'b00, 2'b00, 2'b01, 2'b00, 2'b00, 2'b00, 2'b00, 2'b01, 2'b11, 2'b11, 2'b01, 2'b00, 2'b00, 2'b10, 2'b01, 2'b01, 2'b00, 2'b01, 2'b11, 2'b11, 2'b00, 2'b11, 2'b01, 2'b11, 2'b11, 2'b00, 2'b01 },
		'{ 2'b01, 2'b01, 2'b11, 2'b11, 2'b01, 2'b11, 2'b11, 2'b00, 2'b01, 2'b00, 2'b11, 2'b11, 2'b00, 2'b11, 2'b01, 2'b11, 2'b00, 2'b11, 2'b00, 2'b00, 2'b11, 2'b11, 2'b00, 2'b01, 2'b11, 2'b01, 2'b00, 2'b00, 2'b00, 2'b01, 2'b01, 2'b10, 2'b11, 2'b01, 2'b00, 2'b01, 2'b00, 2'b01, 2'b00, 2'b10, 2'b01, 2'b00, 2'b00, 2'b00, 2'b01, 2'b11, 2'b00, 2'b00, 2'b00, 2'b01, 2'b10, 2'b11, 2'b11, 2'b01, 2'b00, 2'b00, 2'b00, 2'b01, 2'b00, 2'b00, 2'b00, 2'b11, 2'b01, 2'b10 },
		'{ 2'b01, 2'b01, 2'b01, 2'b11, 2'b11, 2'b01, 2'b01, 2'b11, 2'b00, 2'b01, 2'b11, 2'b01, 2'b10, 2'b01, 2'b11, 2'b10, 2'b11, 2'b00, 2'b00, 2'b00, 2'b00, 2'b11, 2'b00, 2'b11, 2'b11, 2'b00, 2'b01, 2'b00, 2'b00, 2'b11, 2'b01, 2'b01, 2'b01, 2'b00, 2'b00, 2'b01, 2'b11, 2'b00, 2'b00, 2'b00, 2'b11, 2'b11, 2'b00, 2'b01, 2'b10, 2'b11, 2'b00, 2'b11, 2'b00, 2'b00, 2'b00, 2'b01, 2'b01, 2'b00, 2'b00, 2'b00, 2'b00, 2'b11, 2'b00, 2'b01, 2'b11, 2'b00, 2'b00, 2'b00 },
		'{ 2'b01, 2'b01, 2'b00, 2'b10, 2'b01, 2'b00, 2'b00, 2'b00, 2'b00, 2'b00, 2'b01, 2'b01, 2'b01, 2'b00, 2'b01, 2'b00, 2'b00, 2'b10, 2'b00, 2'b11, 2'b00, 2'b01, 2'b01, 2'b00, 2'b01, 2'b01, 2'b11, 2'b01, 2'b11, 2'b01, 2'b01, 2'b10, 2'b10, 2'b01, 2'b00, 2'b00, 2'b00, 2'b10, 2'b00, 2'b00, 2'b11, 2'b11, 2'b11, 2'b01, 2'b11, 2'b01, 2'b11, 2'b11, 2'b11, 2'b00, 2'b00, 2'b11, 2'b00, 2'b10, 2'b00, 2'b00, 2'b11, 2'b10, 2'b01, 2'b00, 2'b10, 2'b00, 2'b00, 2'b10 },
		'{ 2'b00, 2'b11, 2'b00, 2'b00, 2'b00, 2'b11, 2'b11, 2'b01, 2'b00, 2'b11, 2'b11, 2'b01, 2'b00, 2'b01, 2'b00, 2'b00, 2'b00, 2'b01, 2'b11, 2'b01, 2'b00, 2'b00, 2'b11, 2'b00, 2'b00, 2'b01, 2'b00, 2'b01, 2'b01, 2'b01, 2'b11, 2'b11, 2'b00, 2'b00, 2'b10, 2'b00, 2'b11, 2'b00, 2'b00, 2'b00, 2'b01, 2'b01, 2'b00, 2'b01, 2'b11, 2'b01, 2'b01, 2'b01, 2'b00, 2'b11, 2'b01, 2'b00, 2'b01, 2'b10, 2'b11, 2'b00, 2'b00, 2'b11, 2'b10, 2'b11, 2'b11, 2'b01, 2'b00, 2'b01 },
		'{ 2'b11, 2'b00, 2'b00, 2'b00, 2'b00, 2'b11, 2'b01, 2'b01, 2'b01, 2'b00, 2'b00, 2'b00, 2'b00, 2'b00, 2'b11, 2'b00, 2'b00, 2'b00, 2'b00, 2'b01, 2'b00, 2'b00, 2'b11, 2'b01, 2'b00, 2'b11, 2'b11, 2'b00, 2'b01, 2'b01, 2'b00, 2'b11, 2'b00, 2'b00, 2'b00, 2'b11, 2'b11, 2'b00, 2'b00, 2'b11, 2'b00, 2'b11, 2'b00, 2'b00, 2'b11, 2'b00, 2'b01, 2'b01, 2'b01, 2'b11, 2'b11, 2'b11, 2'b00, 2'b00, 2'b00, 2'b11, 2'b00, 2'b01, 2'b11, 2'b11, 2'b00, 2'b11, 2'b11, 2'b00 },
		'{ 2'b00, 2'b00, 2'b01, 2'b10, 2'b01, 2'b00, 2'b11, 2'b11, 2'b00, 2'b00, 2'b00, 2'b00, 2'b00, 2'b00, 2'b00, 2'b00, 2'b10, 2'b11, 2'b10, 2'b10, 2'b01, 2'b11, 2'b00, 2'b01, 2'b00, 2'b01, 2'b01, 2'b00, 2'b11, 2'b00, 2'b01, 2'b00, 2'b11, 2'b00, 2'b00, 2'b10, 2'b00, 2'b01, 2'b01, 2'b00, 2'b01, 2'b00, 2'b11, 2'b00, 2'b00, 2'b01, 2'b00, 2'b00, 2'b11, 2'b01, 2'b01, 2'b00, 2'b11, 2'b01, 2'b00, 2'b00, 2'b10, 2'b01, 2'b11, 2'b11, 2'b01, 2'b11, 2'b10, 2'b00 },
		'{ 2'b01, 2'b00, 2'b01, 2'b01, 2'b01, 2'b01, 2'b11, 2'b10, 2'b00, 2'b00, 2'b01, 2'b00, 2'b01, 2'b11, 2'b00, 2'b11, 2'b01, 2'b11, 2'b10, 2'b00, 2'b01, 2'b11, 2'b11, 2'b00, 2'b01, 2'b11, 2'b00, 2'b11, 2'b00, 2'b01, 2'b11, 2'b11, 2'b01, 2'b01, 2'b01, 2'b00, 2'b01, 2'b01, 2'b01, 2'b00, 2'b01, 2'b11, 2'b01, 2'b00, 2'b01, 2'b01, 2'b11, 2'b11, 2'b01, 2'b00, 2'b00, 2'b11, 2'b11, 2'b01, 2'b11, 2'b00, 2'b11, 2'b00, 2'b01, 2'b00, 2'b00, 2'b11, 2'b00, 2'b00 },
		'{ 2'b10, 2'b00, 2'b00, 2'b01, 2'b00, 2'b01, 2'b00, 2'b11, 2'b00, 2'b11, 2'b01, 2'b00, 2'b11, 2'b00, 2'b11, 2'b01, 2'b01, 2'b01, 2'b00, 2'b11, 2'b11, 2'b00, 2'b00, 2'b11, 2'b00, 2'b11, 2'b01, 2'b01, 2'b11, 2'b01, 2'b00, 2'b11, 2'b00, 2'b11, 2'b00, 2'b10, 2'b11, 2'b00, 2'b11, 2'b01, 2'b01, 2'b11, 2'b01, 2'b00, 2'b11, 2'b00, 2'b00, 2'b01, 2'b00, 2'b11, 2'b01, 2'b11, 2'b01, 2'b00, 2'b01, 2'b01, 2'b01, 2'b00, 2'b00, 2'b00, 2'b11, 2'b01, 2'b00, 2'b11 },
		'{ 2'b11, 2'b00, 2'b01, 2'b10, 2'b01, 2'b00, 2'b00, 2'b01, 2'b00, 2'b01, 2'b00, 2'b00, 2'b00, 2'b00, 2'b00, 2'b00, 2'b01, 2'b00, 2'b01, 2'b10, 2'b10, 2'b00, 2'b11, 2'b11, 2'b10, 2'b11, 2'b11, 2'b11, 2'b00, 2'b00, 2'b10, 2'b01, 2'b00, 2'b10, 2'b01, 2'b10, 2'b00, 2'b10, 2'b00, 2'b01, 2'b11, 2'b11, 2'b00, 2'b01, 2'b00, 2'b01, 2'b11, 2'b10, 2'b11, 2'b11, 2'b01, 2'b00, 2'b00, 2'b11, 2'b01, 2'b00, 2'b01, 2'b00, 2'b11, 2'b01, 2'b01, 2'b10, 2'b01, 2'b11 },
		'{ 2'b11, 2'b00, 2'b01, 2'b11, 2'b00, 2'b00, 2'b00, 2'b01, 2'b01, 2'b00, 2'b10, 2'b00, 2'b01, 2'b01, 2'b11, 2'b01, 2'b00, 2'b11, 2'b00, 2'b00, 2'b10, 2'b10, 2'b10, 2'b00, 2'b01, 2'b01, 2'b11, 2'b01, 2'b11, 2'b01, 2'b01, 2'b00, 2'b01, 2'b00, 2'b10, 2'b00, 2'b10, 2'b01, 2'b01, 2'b11, 2'b01, 2'b00, 2'b11, 2'b11, 2'b11, 2'b01, 2'b00, 2'b01, 2'b01, 2'b11, 2'b11, 2'b01, 2'b00, 2'b00, 2'b11, 2'b00, 2'b01, 2'b00, 2'b11, 2'b00, 2'b01, 2'b00, 2'b01, 2'b00 },
		'{ 2'b00, 2'b11, 2'b00, 2'b00, 2'b00, 2'b01, 2'b01, 2'b00, 2'b01, 2'b11, 2'b01, 2'b01, 2'b00, 2'b01, 2'b00, 2'b11, 2'b00, 2'b11, 2'b00, 2'b11, 2'b00, 2'b11, 2'b00, 2'b01, 2'b10, 2'b00, 2'b11, 2'b01, 2'b11, 2'b01, 2'b10, 2'b00, 2'b00, 2'b00, 2'b11, 2'b10, 2'b01, 2'b00, 2'b01, 2'b10, 2'b11, 2'b01, 2'b10, 2'b00, 2'b10, 2'b00, 2'b00, 2'b01, 2'b01, 2'b00, 2'b00, 2'b10, 2'b00, 2'b01, 2'b01, 2'b00, 2'b00, 2'b11, 2'b10, 2'b00, 2'b01, 2'b10, 2'b00, 2'b00 },
		'{ 2'b00, 2'b00, 2'b11, 2'b01, 2'b00, 2'b00, 2'b01, 2'b00, 2'b01, 2'b11, 2'b00, 2'b11, 2'b11, 2'b10, 2'b11, 2'b01, 2'b11, 2'b11, 2'b11, 2'b11, 2'b01, 2'b00, 2'b10, 2'b00, 2'b00, 2'b11, 2'b10, 2'b01, 2'b00, 2'b00, 2'b01, 2'b10, 2'b00, 2'b11, 2'b01, 2'b00, 2'b11, 2'b10, 2'b01, 2'b00, 2'b00, 2'b01, 2'b00, 2'b00, 2'b11, 2'b00, 2'b01, 2'b01, 2'b00, 2'b11, 2'b11, 2'b11, 2'b01, 2'b01, 2'b01, 2'b00, 2'b11, 2'b00, 2'b00, 2'b00, 2'b01, 2'b01, 2'b01, 2'b00 },
		'{ 2'b01, 2'b00, 2'b00, 2'b00, 2'b11, 2'b00, 2'b11, 2'b10, 2'b00, 2'b10, 2'b01, 2'b01, 2'b01, 2'b11, 2'b01, 2'b10, 2'b11, 2'b11, 2'b01, 2'b01, 2'b11, 2'b00, 2'b01, 2'b11, 2'b00, 2'b00, 2'b01, 2'b01, 2'b00, 2'b11, 2'b00, 2'b00, 2'b01, 2'b11, 2'b11, 2'b01, 2'b00, 2'b01, 2'b10, 2'b00, 2'b00, 2'b00, 2'b00, 2'b10, 2'b01, 2'b00, 2'b00, 2'b10, 2'b01, 2'b00, 2'b01, 2'b11, 2'b11, 2'b11, 2'b01, 2'b11, 2'b01, 2'b11, 2'b11, 2'b01, 2'b01, 2'b11, 2'b00, 2'b11 },
		'{ 2'b10, 2'b00, 2'b00, 2'b01, 2'b00, 2'b11, 2'b01, 2'b11, 2'b00, 2'b00, 2'b01, 2'b01, 2'b00, 2'b01, 2'b01, 2'b00, 2'b01, 2'b01, 2'b00, 2'b00, 2'b01, 2'b00, 2'b01, 2'b00, 2'b11, 2'b11, 2'b01, 2'b01, 2'b00, 2'b00, 2'b10, 2'b00, 2'b00, 2'b01, 2'b01, 2'b11, 2'b11, 2'b01, 2'b10, 2'b00, 2'b01, 2'b11, 2'b11, 2'b01, 2'b11, 2'b00, 2'b01, 2'b11, 2'b01, 2'b01, 2'b11, 2'b00, 2'b11, 2'b00, 2'b01, 2'b00, 2'b00, 2'b10, 2'b01, 2'b01, 2'b00, 2'b10, 2'b10, 2'b00 },
		'{ 2'b01, 2'b11, 2'b11, 2'b00, 2'b01, 2'b00, 2'b00, 2'b11, 2'b00, 2'b11, 2'b00, 2'b11, 2'b01, 2'b00, 2'b00, 2'b11, 2'b00, 2'b01, 2'b01, 2'b00, 2'b10, 2'b01, 2'b01, 2'b11, 2'b00, 2'b01, 2'b01, 2'b10, 2'b01, 2'b01, 2'b11, 2'b00, 2'b00, 2'b00, 2'b00, 2'b01, 2'b00, 2'b11, 2'b11, 2'b11, 2'b11, 2'b00, 2'b00, 2'b11, 2'b11, 2'b00, 2'b11, 2'b00, 2'b00, 2'b00, 2'b11, 2'b10, 2'b00, 2'b01, 2'b00, 2'b01, 2'b00, 2'b11, 2'b01, 2'b11, 2'b00, 2'b01, 2'b00, 2'b11 },
		'{ 2'b10, 2'b01, 2'b01, 2'b11, 2'b11, 2'b01, 2'b11, 2'b11, 2'b11, 2'b00, 2'b01, 2'b01, 2'b10, 2'b01, 2'b00, 2'b11, 2'b01, 2'b01, 2'b10, 2'b00, 2'b00, 2'b01, 2'b00, 2'b00, 2'b11, 2'b00, 2'b00, 2'b01, 2'b11, 2'b00, 2'b11, 2'b00, 2'b01, 2'b00, 2'b11, 2'b01, 2'b11, 2'b11, 2'b01, 2'b00, 2'b00, 2'b11, 2'b01, 2'b01, 2'b11, 2'b01, 2'b11, 2'b10, 2'b00, 2'b11, 2'b00, 2'b10, 2'b00, 2'b11, 2'b01, 2'b11, 2'b01, 2'b11, 2'b11, 2'b10, 2'b01, 2'b11, 2'b01, 2'b00 },
		'{ 2'b11, 2'b11, 2'b11, 2'b01, 2'b00, 2'b10, 2'b00, 2'b10, 2'b00, 2'b01, 2'b11, 2'b00, 2'b01, 2'b00, 2'b01, 2'b01, 2'b11, 2'b01, 2'b01, 2'b00, 2'b01, 2'b00, 2'b01, 2'b00, 2'b01, 2'b01, 2'b00, 2'b11, 2'b00, 2'b00, 2'b01, 2'b01, 2'b00, 2'b01, 2'b01, 2'b11, 2'b11, 2'b01, 2'b00, 2'b11, 2'b01, 2'b01, 2'b00, 2'b11, 2'b01, 2'b01, 2'b00, 2'b11, 2'b11, 2'b10, 2'b01, 2'b10, 2'b01, 2'b00, 2'b11, 2'b01, 2'b00, 2'b01, 2'b10, 2'b11, 2'b01, 2'b01, 2'b00, 2'b11 },
		'{ 2'b10, 2'b01, 2'b01, 2'b01, 2'b11, 2'b00, 2'b01, 2'b01, 2'b00, 2'b00, 2'b01, 2'b11, 2'b01, 2'b01, 2'b01, 2'b00, 2'b00, 2'b11, 2'b10, 2'b01, 2'b00, 2'b00, 2'b00, 2'b10, 2'b00, 2'b00, 2'b10, 2'b01, 2'b01, 2'b11, 2'b00, 2'b00, 2'b00, 2'b00, 2'b01, 2'b01, 2'b00, 2'b01, 2'b00, 2'b00, 2'b00, 2'b00, 2'b01, 2'b01, 2'b01, 2'b00, 2'b00, 2'b11, 2'b10, 2'b00, 2'b00, 2'b00, 2'b00, 2'b01, 2'b01, 2'b00, 2'b00, 2'b11, 2'b11, 2'b01, 2'b00, 2'b00, 2'b01, 2'b00 },
		'{ 2'b11, 2'b10, 2'b01, 2'b00, 2'b01, 2'b00, 2'b00, 2'b00, 2'b01, 2'b11, 2'b11, 2'b00, 2'b01, 2'b01, 2'b01, 2'b01, 2'b11, 2'b11, 2'b11, 2'b00, 2'b00, 2'b10, 2'b01, 2'b00, 2'b01, 2'b01, 2'b00, 2'b11, 2'b00, 2'b11, 2'b11, 2'b11, 2'b00, 2'b00, 2'b01, 2'b00, 2'b00, 2'b00, 2'b01, 2'b00, 2'b11, 2'b10, 2'b11, 2'b11, 2'b01, 2'b00, 2'b01, 2'b01, 2'b01, 2'b01, 2'b10, 2'b11, 2'b00, 2'b11, 2'b00, 2'b01, 2'b00, 2'b00, 2'b10, 2'b01, 2'b01, 2'b01, 2'b11, 2'b00 },
		'{ 2'b01, 2'b11, 2'b10, 2'b11, 2'b00, 2'b01, 2'b00, 2'b11, 2'b00, 2'b11, 2'b00, 2'b01, 2'b01, 2'b11, 2'b00, 2'b01, 2'b11, 2'b00, 2'b11, 2'b11, 2'b01, 2'b10, 2'b01, 2'b01, 2'b00, 2'b11, 2'b00, 2'b00, 2'b01, 2'b01, 2'b01, 2'b00, 2'b11, 2'b01, 2'b00, 2'b00, 2'b00, 2'b00, 2'b11, 2'b00, 2'b11, 2'b11, 2'b11, 2'b11, 2'b10, 2'b01, 2'b01, 2'b11, 2'b01, 2'b00, 2'b01, 2'b01, 2'b11, 2'b00, 2'b00, 2'b01, 2'b01, 2'b00, 2'b01, 2'b11, 2'b01, 2'b11, 2'b11, 2'b10 },
		'{ 2'b01, 2'b01, 2'b10, 2'b00, 2'b00, 2'b00, 2'b10, 2'b10, 2'b11, 2'b00, 2'b00, 2'b00, 2'b01, 2'b00, 2'b00, 2'b00, 2'b01, 2'b00, 2'b01, 2'b01, 2'b00, 2'b01, 2'b00, 2'b00, 2'b00, 2'b11, 2'b00, 2'b11, 2'b01, 2'b01, 2'b10, 2'b10, 2'b01, 2'b00, 2'b11, 2'b01, 2'b11, 2'b00, 2'b10, 2'b11, 2'b01, 2'b11, 2'b00, 2'b01, 2'b11, 2'b11, 2'b11, 2'b00, 2'b11, 2'b00, 2'b01, 2'b00, 2'b00, 2'b01, 2'b01, 2'b01, 2'b11, 2'b00, 2'b00, 2'b11, 2'b00, 2'b01, 2'b00, 2'b00 },
		'{ 2'b00, 2'b11, 2'b01, 2'b00, 2'b00, 2'b00, 2'b01, 2'b01, 2'b11, 2'b01, 2'b00, 2'b01, 2'b01, 2'b01, 2'b10, 2'b01, 2'b00, 2'b10, 2'b10, 2'b01, 2'b11, 2'b01, 2'b00, 2'b01, 2'b00, 2'b01, 2'b11, 2'b00, 2'b00, 2'b11, 2'b00, 2'b10, 2'b01, 2'b00, 2'b01, 2'b11, 2'b11, 2'b10, 2'b00, 2'b01, 2'b11, 2'b11, 2'b00, 2'b00, 2'b00, 2'b01, 2'b01, 2'b01, 2'b00, 2'b11, 2'b01, 2'b00, 2'b00, 2'b00, 2'b00, 2'b11, 2'b11, 2'b00, 2'b11, 2'b00, 2'b01, 2'b11, 2'b00, 2'b01 },
		'{ 2'b00, 2'b01, 2'b11, 2'b11, 2'b00, 2'b11, 2'b00, 2'b01, 2'b00, 2'b01, 2'b11, 2'b10, 2'b10, 2'b00, 2'b11, 2'b11, 2'b00, 2'b11, 2'b10, 2'b11, 2'b01, 2'b00, 2'b01, 2'b00, 2'b11, 2'b00, 2'b11, 2'b00, 2'b00, 2'b11, 2'b11, 2'b01, 2'b01, 2'b00, 2'b00, 2'b11, 2'b00, 2'b01, 2'b00, 2'b11, 2'b01, 2'b00, 2'b00, 2'b11, 2'b00, 2'b10, 2'b01, 2'b11, 2'b11, 2'b00, 2'b01, 2'b11, 2'b11, 2'b00, 2'b11, 2'b00, 2'b01, 2'b01, 2'b00, 2'b00, 2'b00, 2'b00, 2'b01, 2'b11 },
		'{ 2'b00, 2'b00, 2'b01, 2'b01, 2'b01, 2'b00, 2'b00, 2'b00, 2'b00, 2'b00, 2'b10, 2'b00, 2'b01, 2'b01, 2'b01, 2'b00, 2'b00, 2'b11, 2'b01, 2'b00, 2'b01, 2'b00, 2'b01, 2'b01, 2'b11, 2'b01, 2'b01, 2'b11, 2'b00, 2'b01, 2'b00, 2'b11, 2'b01, 2'b00, 2'b00, 2'b00, 2'b01, 2'b00, 2'b10, 2'b01, 2'b10, 2'b00, 2'b00, 2'b11, 2'b00, 2'b01, 2'b11, 2'b00, 2'b11, 2'b11, 2'b01, 2'b01, 2'b11, 2'b01, 2'b01, 2'b10, 2'b00, 2'b11, 2'b00, 2'b00, 2'b01, 2'b01, 2'b11, 2'b01 },
		'{ 2'b00, 2'b11, 2'b01, 2'b11, 2'b00, 2'b00, 2'b11, 2'b00, 2'b11, 2'b01, 2'b01, 2'b01, 2'b00, 2'b00, 2'b11, 2'b01, 2'b11, 2'b11, 2'b00, 2'b11, 2'b00, 2'b01, 2'b01, 2'b00, 2'b00, 2'b00, 2'b01, 2'b00, 2'b01, 2'b11, 2'b11, 2'b01, 2'b00, 2'b10, 2'b00, 2'b01, 2'b00, 2'b00, 2'b11, 2'b01, 2'b00, 2'b10, 2'b00, 2'b01, 2'b01, 2'b01, 2'b11, 2'b00, 2'b01, 2'b00, 2'b01, 2'b00, 2'b00, 2'b01, 2'b01, 2'b00, 2'b01, 2'b00, 2'b01, 2'b00, 2'b01, 2'b01, 2'b01, 2'b00 },
		'{ 2'b01, 2'b00, 2'b01, 2'b01, 2'b11, 2'b00, 2'b01, 2'b11, 2'b01, 2'b11, 2'b00, 2'b10, 2'b11, 2'b11, 2'b01, 2'b00, 2'b01, 2'b01, 2'b11, 2'b00, 2'b11, 2'b01, 2'b00, 2'b01, 2'b00, 2'b00, 2'b01, 2'b01, 2'b01, 2'b11, 2'b01, 2'b10, 2'b01, 2'b11, 2'b01, 2'b00, 2'b11, 2'b00, 2'b01, 2'b01, 2'b00, 2'b11, 2'b01, 2'b00, 2'b00, 2'b11, 2'b11, 2'b01, 2'b00, 2'b00, 2'b10, 2'b00, 2'b11, 2'b00, 2'b01, 2'b10, 2'b10, 2'b01, 2'b00, 2'b00, 2'b11, 2'b11, 2'b01, 2'b11 },
		'{ 2'b00, 2'b00, 2'b00, 2'b00, 2'b00, 2'b01, 2'b10, 2'b11, 2'b11, 2'b01, 2'b00, 2'b01, 2'b00, 2'b00, 2'b00, 2'b00, 2'b00, 2'b00, 2'b01, 2'b01, 2'b11, 2'b00, 2'b00, 2'b00, 2'b11, 2'b00, 2'b11, 2'b00, 2'b11, 2'b01, 2'b01, 2'b01, 2'b10, 2'b11, 2'b11, 2'b00, 2'b00, 2'b00, 2'b01, 2'b00, 2'b10, 2'b00, 2'b11, 2'b00, 2'b00, 2'b11, 2'b00, 2'b11, 2'b11, 2'b00, 2'b11, 2'b00, 2'b00, 2'b00, 2'b01, 2'b11, 2'b00, 2'b00, 2'b11, 2'b00, 2'b00, 2'b01, 2'b00, 2'b00 },
		'{ 2'b01, 2'b00, 2'b11, 2'b11, 2'b11, 2'b01, 2'b00, 2'b01, 2'b10, 2'b01, 2'b11, 2'b11, 2'b01, 2'b10, 2'b11, 2'b01, 2'b01, 2'b11, 2'b00, 2'b11, 2'b01, 2'b11, 2'b00, 2'b10, 2'b01, 2'b01, 2'b00, 2'b00, 2'b11, 2'b01, 2'b00, 2'b00, 2'b11, 2'b11, 2'b10, 2'b00, 2'b10, 2'b10, 2'b01, 2'b01, 2'b10, 2'b00, 2'b11, 2'b11, 2'b01, 2'b00, 2'b00, 2'b00, 2'b11, 2'b11, 2'b00, 2'b01, 2'b00, 2'b11, 2'b11, 2'b00, 2'b01, 2'b00, 2'b11, 2'b00, 2'b01, 2'b00, 2'b01, 2'b01 },
		'{ 2'b00, 2'b00, 2'b01, 2'b01, 2'b01, 2'b00, 2'b01, 2'b00, 2'b01, 2'b01, 2'b00, 2'b00, 2'b11, 2'b01, 2'b11, 2'b01, 2'b10, 2'b01, 2'b10, 2'b00, 2'b11, 2'b00, 2'b00, 2'b10, 2'b10, 2'b00, 2'b11, 2'b01, 2'b00, 2'b00, 2'b01, 2'b00, 2'b00, 2'b00, 2'b00, 2'b00, 2'b01, 2'b01, 2'b00, 2'b11, 2'b01, 2'b00, 2'b11, 2'b00, 2'b00, 2'b11, 2'b11, 2'b01, 2'b00, 2'b00, 2'b10, 2'b00, 2'b11, 2'b00, 2'b00, 2'b11, 2'b11, 2'b01, 2'b11, 2'b00, 2'b00, 2'b01, 2'b11, 2'b01 },
		'{ 2'b00, 2'b01, 2'b11, 2'b00, 2'b10, 2'b00, 2'b11, 2'b10, 2'b10, 2'b00, 2'b00, 2'b01, 2'b11, 2'b00, 2'b01, 2'b01, 2'b00, 2'b01, 2'b00, 2'b00, 2'b10, 2'b00, 2'b11, 2'b11, 2'b01, 2'b01, 2'b00, 2'b11, 2'b01, 2'b01, 2'b10, 2'b00, 2'b11, 2'b00, 2'b00, 2'b00, 2'b11, 2'b00, 2'b11, 2'b10, 2'b11, 2'b00, 2'b00, 2'b00, 2'b00, 2'b11, 2'b00, 2'b00, 2'b10, 2'b11, 2'b11, 2'b00, 2'b00, 2'b00, 2'b01, 2'b00, 2'b01, 2'b11, 2'b00, 2'b11, 2'b01, 2'b00, 2'b11, 2'b01 },
		'{ 2'b01, 2'b00, 2'b11, 2'b00, 2'b10, 2'b01, 2'b01, 2'b01, 2'b01, 2'b10, 2'b00, 2'b10, 2'b11, 2'b00, 2'b00, 2'b00, 2'b00, 2'b10, 2'b00, 2'b01, 2'b11, 2'b00, 2'b00, 2'b11, 2'b01, 2'b11, 2'b11, 2'b11, 2'b00, 2'b01, 2'b00, 2'b00, 2'b11, 2'b00, 2'b01, 2'b01, 2'b01, 2'b10, 2'b11, 2'b00, 2'b01, 2'b01, 2'b01, 2'b11, 2'b01, 2'b01, 2'b00, 2'b01, 2'b00, 2'b01, 2'b01, 2'b11, 2'b01, 2'b11, 2'b01, 2'b01, 2'b11, 2'b11, 2'b00, 2'b00, 2'b00, 2'b11, 2'b01, 2'b00 },
		'{ 2'b00, 2'b01, 2'b01, 2'b00, 2'b00, 2'b00, 2'b01, 2'b01, 2'b00, 2'b11, 2'b00, 2'b01, 2'b01, 2'b01, 2'b11, 2'b01, 2'b01, 2'b01, 2'b11, 2'b11, 2'b00, 2'b01, 2'b01, 2'b00, 2'b11, 2'b10, 2'b01, 2'b11, 2'b01, 2'b00, 2'b11, 2'b11, 2'b10, 2'b10, 2'b10, 2'b00, 2'b00, 2'b00, 2'b11, 2'b00, 2'b10, 2'b11, 2'b11, 2'b01, 2'b11, 2'b11, 2'b11, 2'b00, 2'b11, 2'b01, 2'b00, 2'b01, 2'b00, 2'b01, 2'b01, 2'b01, 2'b01, 2'b00, 2'b01, 2'b01, 2'b11, 2'b00, 2'b01, 2'b11 },
		'{ 2'b00, 2'b00, 2'b11, 2'b11, 2'b01, 2'b11, 2'b11, 2'b11, 2'b10, 2'b01, 2'b00, 2'b01, 2'b00, 2'b10, 2'b01, 2'b11, 2'b00, 2'b11, 2'b11, 2'b00, 2'b11, 2'b00, 2'b01, 2'b10, 2'b11, 2'b11, 2'b01, 2'b01, 2'b10, 2'b01, 2'b00, 2'b11, 2'b11, 2'b01, 2'b00, 2'b11, 2'b01, 2'b00, 2'b11, 2'b11, 2'b11, 2'b11, 2'b00, 2'b00, 2'b01, 2'b11, 2'b00, 2'b11, 2'b00, 2'b11, 2'b10, 2'b01, 2'b01, 2'b00, 2'b11, 2'b11, 2'b11, 2'b00, 2'b00, 2'b11, 2'b00, 2'b00, 2'b00, 2'b01 },
		'{ 2'b00, 2'b01, 2'b10, 2'b01, 2'b00, 2'b11, 2'b00, 2'b00, 2'b00, 2'b00, 2'b00, 2'b10, 2'b01, 2'b00, 2'b11, 2'b00, 2'b01, 2'b01, 2'b00, 2'b01, 2'b11, 2'b01, 2'b00, 2'b01, 2'b11, 2'b10, 2'b01, 2'b01, 2'b00, 2'b01, 2'b01, 2'b00, 2'b11, 2'b00, 2'b00, 2'b01, 2'b10, 2'b00, 2'b10, 2'b01, 2'b00, 2'b01, 2'b10, 2'b10, 2'b11, 2'b01, 2'b10, 2'b01, 2'b00, 2'b00, 2'b10, 2'b10, 2'b11, 2'b11, 2'b00, 2'b00, 2'b01, 2'b01, 2'b00, 2'b00, 2'b00, 2'b11, 2'b00, 2'b00 },
		'{ 2'b00, 2'b01, 2'b01, 2'b00, 2'b00, 2'b00, 2'b11, 2'b11, 2'b01, 2'b01, 2'b01, 2'b11, 2'b01, 2'b11, 2'b01, 2'b00, 2'b00, 2'b11, 2'b01, 2'b11, 2'b01, 2'b01, 2'b11, 2'b00, 2'b00, 2'b11, 2'b00, 2'b01, 2'b01, 2'b00, 2'b01, 2'b01, 2'b11, 2'b00, 2'b00, 2'b00, 2'b00, 2'b11, 2'b01, 2'b10, 2'b01, 2'b01, 2'b11, 2'b01, 2'b11, 2'b00, 2'b00, 2'b00, 2'b00, 2'b11, 2'b00, 2'b01, 2'b00, 2'b01, 2'b00, 2'b11, 2'b00, 2'b00, 2'b01, 2'b00, 2'b00, 2'b11, 2'b01, 2'b00 },
		'{ 2'b11, 2'b00, 2'b01, 2'b00, 2'b11, 2'b01, 2'b11, 2'b11, 2'b11, 2'b01, 2'b01, 2'b11, 2'b01, 2'b00, 2'b01, 2'b00, 2'b01, 2'b11, 2'b01, 2'b01, 2'b00, 2'b11, 2'b01, 2'b01, 2'b01, 2'b00, 2'b11, 2'b01, 2'b00, 2'b01, 2'b01, 2'b01, 2'b01, 2'b00, 2'b01, 2'b11, 2'b11, 2'b10, 2'b10, 2'b00, 2'b01, 2'b11, 2'b01, 2'b00, 2'b00, 2'b00, 2'b01, 2'b11, 2'b01, 2'b00, 2'b01, 2'b01, 2'b01, 2'b10, 2'b00, 2'b11, 2'b11, 2'b00, 2'b00, 2'b01, 2'b00, 2'b01, 2'b01, 2'b01 },
		'{ 2'b01, 2'b01, 2'b01, 2'b00, 2'b00, 2'b01, 2'b00, 2'b10, 2'b00, 2'b00, 2'b00, 2'b01, 2'b00, 2'b01, 2'b01, 2'b01, 2'b01, 2'b00, 2'b00, 2'b01, 2'b01, 2'b11, 2'b10, 2'b00, 2'b01, 2'b11, 2'b01, 2'b01, 2'b00, 2'b10, 2'b00, 2'b10, 2'b00, 2'b01, 2'b01, 2'b00, 2'b11, 2'b00, 2'b11, 2'b10, 2'b01, 2'b00, 2'b11, 2'b01, 2'b01, 2'b00, 2'b01, 2'b10, 2'b01, 2'b11, 2'b01, 2'b00, 2'b01, 2'b00, 2'b00, 2'b11, 2'b01, 2'b01, 2'b01, 2'b01, 2'b11, 2'b00, 2'b00, 2'b11 },
		'{ 2'b11, 2'b01, 2'b00, 2'b01, 2'b00, 2'b00, 2'b00, 2'b11, 2'b01, 2'b00, 2'b00, 2'b00, 2'b00, 2'b11, 2'b11, 2'b00, 2'b11, 2'b00, 2'b11, 2'b00, 2'b01, 2'b01, 2'b01, 2'b01, 2'b11, 2'b01, 2'b00, 2'b11, 2'b00, 2'b00, 2'b01, 2'b00, 2'b00, 2'b01, 2'b00, 2'b00, 2'b11, 2'b00, 2'b00, 2'b00, 2'b00, 2'b11, 2'b00, 2'b10, 2'b11, 2'b11, 2'b11, 2'b10, 2'b01, 2'b00, 2'b01, 2'b01, 2'b01, 2'b00, 2'b00, 2'b11, 2'b00, 2'b01, 2'b00, 2'b00, 2'b01, 2'b10, 2'b11, 2'b00 },
		'{ 2'b00, 2'b01, 2'b00, 2'b00, 2'b01, 2'b01, 2'b01, 2'b11, 2'b11, 2'b00, 2'b00, 2'b01, 2'b10, 2'b00, 2'b01, 2'b00, 2'b00, 2'b00, 2'b01, 2'b01, 2'b01, 2'b00, 2'b00, 2'b11, 2'b01, 2'b00, 2'b01, 2'b00, 2'b00, 2'b01, 2'b01, 2'b11, 2'b01, 2'b11, 2'b11, 2'b01, 2'b00, 2'b00, 2'b00, 2'b00, 2'b00, 2'b00, 2'b00, 2'b01, 2'b11, 2'b01, 2'b01, 2'b00, 2'b00, 2'b01, 2'b00, 2'b01, 2'b00, 2'b00, 2'b00, 2'b11, 2'b00, 2'b11, 2'b10, 2'b01, 2'b01, 2'b01, 2'b00, 2'b01 },
		'{ 2'b11, 2'b11, 2'b01, 2'b00, 2'b01, 2'b00, 2'b00, 2'b10, 2'b00, 2'b00, 2'b11, 2'b00, 2'b01, 2'b10, 2'b00, 2'b00, 2'b01, 2'b00, 2'b01, 2'b01, 2'b01, 2'b01, 2'b00, 2'b00, 2'b11, 2'b01, 2'b01, 2'b00, 2'b00, 2'b00, 2'b11, 2'b11, 2'b11, 2'b10, 2'b11, 2'b10, 2'b00, 2'b00, 2'b01, 2'b11, 2'b10, 2'b00, 2'b11, 2'b00, 2'b01, 2'b01, 2'b00, 2'b11, 2'b00, 2'b00, 2'b00, 2'b11, 2'b00, 2'b11, 2'b11, 2'b01, 2'b00, 2'b00, 2'b11, 2'b10, 2'b11, 2'b11, 2'b11, 2'b01 },
		'{ 2'b01, 2'b11, 2'b11, 2'b00, 2'b01, 2'b00, 2'b11, 2'b11, 2'b00, 2'b11, 2'b01, 2'b01, 2'b11, 2'b00, 2'b00, 2'b00, 2'b01, 2'b01, 2'b00, 2'b00, 2'b11, 2'b11, 2'b00, 2'b00, 2'b01, 2'b00, 2'b01, 2'b01, 2'b00, 2'b00, 2'b11, 2'b00, 2'b11, 2'b00, 2'b00, 2'b11, 2'b10, 2'b01, 2'b00, 2'b01, 2'b11, 2'b01, 2'b00, 2'b00, 2'b00, 2'b01, 2'b00, 2'b10, 2'b11, 2'b01, 2'b00, 2'b11, 2'b10, 2'b11, 2'b00, 2'b00, 2'b00, 2'b01, 2'b01, 2'b00, 2'b01, 2'b01, 2'b11, 2'b01 },
		'{ 2'b10, 2'b11, 2'b01, 2'b00, 2'b00, 2'b11, 2'b00, 2'b00, 2'b11, 2'b00, 2'b11, 2'b00, 2'b10, 2'b00, 2'b01, 2'b01, 2'b00, 2'b00, 2'b01, 2'b11, 2'b11, 2'b00, 2'b01, 2'b01, 2'b10, 2'b10, 2'b11, 2'b11, 2'b01, 2'b01, 2'b00, 2'b01, 2'b01, 2'b11, 2'b11, 2'b10, 2'b00, 2'b00, 2'b01, 2'b00, 2'b11, 2'b01, 2'b00, 2'b11, 2'b11, 2'b01, 2'b01, 2'b11, 2'b00, 2'b00, 2'b11, 2'b00, 2'b11, 2'b01, 2'b00, 2'b11, 2'b01, 2'b11, 2'b01, 2'b00, 2'b00, 2'b00, 2'b01, 2'b00 },
		'{ 2'b01, 2'b00, 2'b00, 2'b00, 2'b11, 2'b01, 2'b00, 2'b11, 2'b10, 2'b00, 2'b01, 2'b11, 2'b00, 2'b00, 2'b01, 2'b11, 2'b00, 2'b11, 2'b01, 2'b11, 2'b11, 2'b00, 2'b00, 2'b01, 2'b11, 2'b11, 2'b11, 2'b11, 2'b00, 2'b00, 2'b01, 2'b00, 2'b01, 2'b00, 2'b11, 2'b11, 2'b01, 2'b01, 2'b10, 2'b10, 2'b01, 2'b00, 2'b11, 2'b11, 2'b00, 2'b11, 2'b00, 2'b00, 2'b10, 2'b01, 2'b11, 2'b00, 2'b11, 2'b01, 2'b00, 2'b00, 2'b01, 2'b01, 2'b00, 2'b00, 2'b01, 2'b11, 2'b11, 2'b01 },
		'{ 2'b00, 2'b00, 2'b00, 2'b00, 2'b11, 2'b11, 2'b00, 2'b00, 2'b01, 2'b00, 2'b11, 2'b01, 2'b10, 2'b11, 2'b01, 2'b11, 2'b00, 2'b11, 2'b10, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b00, 2'b00, 2'b10, 2'b00, 2'b00, 2'b00, 2'b00, 2'b01, 2'b11, 2'b10, 2'b11, 2'b01, 2'b00, 2'b11, 2'b00, 2'b11, 2'b01, 2'b01, 2'b11, 2'b00, 2'b01, 2'b11, 2'b01, 2'b11, 2'b00, 2'b11, 2'b01, 2'b00, 2'b00, 2'b00, 2'b11, 2'b00, 2'b00, 2'b01, 2'b00, 2'b00, 2'b10, 2'b00, 2'b00, 2'b11 },
		'{ 2'b00, 2'b11, 2'b01, 2'b11, 2'b01, 2'b11, 2'b00, 2'b01, 2'b00, 2'b10, 2'b01, 2'b00, 2'b01, 2'b00, 2'b11, 2'b00, 2'b10, 2'b11, 2'b10, 2'b11, 2'b01, 2'b01, 2'b11, 2'b10, 2'b01, 2'b00, 2'b01, 2'b11, 2'b00, 2'b00, 2'b00, 2'b01, 2'b00, 2'b11, 2'b00, 2'b00, 2'b00, 2'b01, 2'b10, 2'b00, 2'b00, 2'b01, 2'b01, 2'b01, 2'b01, 2'b00, 2'b11, 2'b00, 2'b11, 2'b01, 2'b01, 2'b00, 2'b00, 2'b11, 2'b11, 2'b01, 2'b01, 2'b00, 2'b11, 2'b00, 2'b01, 2'b00, 2'b11, 2'b00 },
		'{ 2'b11, 2'b00, 2'b01, 2'b00, 2'b00, 2'b00, 2'b00, 2'b11, 2'b11, 2'b11, 2'b00, 2'b00, 2'b11, 2'b10, 2'b00, 2'b00, 2'b00, 2'b00, 2'b10, 2'b01, 2'b01, 2'b01, 2'b00, 2'b00, 2'b01, 2'b01, 2'b01, 2'b11, 2'b00, 2'b11, 2'b11, 2'b01, 2'b00, 2'b01, 2'b00, 2'b11, 2'b00, 2'b11, 2'b00, 2'b10, 2'b00, 2'b00, 2'b00, 2'b01, 2'b01, 2'b11, 2'b00, 2'b00, 2'b00, 2'b01, 2'b00, 2'b01, 2'b00, 2'b00, 2'b01, 2'b10, 2'b01, 2'b01, 2'b10, 2'b01, 2'b01, 2'b11, 2'b01, 2'b00 },
		'{ 2'b01, 2'b01, 2'b01, 2'b00, 2'b11, 2'b01, 2'b00, 2'b00, 2'b00, 2'b00, 2'b00, 2'b01, 2'b11, 2'b00, 2'b10, 2'b01, 2'b10, 2'b00, 2'b11, 2'b11, 2'b00, 2'b11, 2'b11, 2'b00, 2'b11, 2'b00, 2'b11, 2'b10, 2'b00, 2'b00, 2'b11, 2'b01, 2'b00, 2'b11, 2'b11, 2'b00, 2'b00, 2'b10, 2'b11, 2'b11, 2'b01, 2'b01, 2'b01, 2'b11, 2'b01, 2'b01, 2'b11, 2'b01, 2'b01, 2'b01, 2'b11, 2'b01, 2'b11, 2'b11, 2'b01, 2'b01, 2'b11, 2'b11, 2'b01, 2'b10, 2'b11, 2'b00, 2'b00, 2'b00 },
		'{ 2'b00, 2'b11, 2'b01, 2'b01, 2'b01, 2'b10, 2'b11, 2'b11, 2'b11, 2'b11, 2'b00, 2'b11, 2'b10, 2'b00, 2'b11, 2'b00, 2'b00, 2'b00, 2'b01, 2'b01, 2'b01, 2'b01, 2'b11, 2'b10, 2'b01, 2'b11, 2'b00, 2'b00, 2'b11, 2'b00, 2'b11, 2'b00, 2'b00, 2'b11, 2'b01, 2'b01, 2'b00, 2'b00, 2'b00, 2'b00, 2'b00, 2'b11, 2'b00, 2'b00, 2'b00, 2'b01, 2'b11, 2'b01, 2'b00, 2'b11, 2'b01, 2'b01, 2'b00, 2'b10, 2'b10, 2'b11, 2'b00, 2'b01, 2'b00, 2'b00, 2'b01, 2'b10, 2'b11, 2'b00 },
		'{ 2'b11, 2'b00, 2'b01, 2'b00, 2'b11, 2'b01, 2'b01, 2'b01, 2'b00, 2'b11, 2'b11, 2'b01, 2'b01, 2'b11, 2'b00, 2'b11, 2'b11, 2'b00, 2'b11, 2'b00, 2'b01, 2'b01, 2'b10, 2'b00, 2'b11, 2'b00, 2'b01, 2'b00, 2'b11, 2'b11, 2'b10, 2'b00, 2'b00, 2'b01, 2'b00, 2'b00, 2'b01, 2'b11, 2'b11, 2'b00, 2'b11, 2'b00, 2'b00, 2'b01, 2'b01, 2'b11, 2'b11, 2'b10, 2'b01, 2'b11, 2'b01, 2'b01, 2'b11, 2'b01, 2'b01, 2'b11, 2'b01, 2'b10, 2'b00, 2'b01, 2'b01, 2'b00, 2'b00, 2'b01 },
		'{ 2'b00, 2'b00, 2'b00, 2'b11, 2'b11, 2'b00, 2'b00, 2'b01, 2'b11, 2'b00, 2'b00, 2'b00, 2'b11, 2'b00, 2'b01, 2'b11, 2'b01, 2'b11, 2'b01, 2'b01, 2'b01, 2'b00, 2'b01, 2'b00, 2'b00, 2'b01, 2'b01, 2'b00, 2'b00, 2'b00, 2'b01, 2'b00, 2'b11, 2'b00, 2'b00, 2'b00, 2'b00, 2'b01, 2'b10, 2'b00, 2'b00, 2'b00, 2'b00, 2'b11, 2'b01, 2'b01, 2'b00, 2'b11, 2'b10, 2'b01, 2'b10, 2'b01, 2'b01, 2'b11, 2'b00, 2'b00, 2'b00, 2'b11, 2'b00, 2'b11, 2'b10, 2'b00, 2'b11, 2'b11 },
		'{ 2'b00, 2'b00, 2'b01, 2'b11, 2'b10, 2'b01, 2'b01, 2'b10, 2'b00, 2'b00, 2'b11, 2'b11, 2'b01, 2'b11, 2'b11, 2'b00, 2'b10, 2'b00, 2'b01, 2'b00, 2'b01, 2'b01, 2'b00, 2'b00, 2'b01, 2'b01, 2'b10, 2'b00, 2'b11, 2'b00, 2'b11, 2'b01, 2'b00, 2'b11, 2'b00, 2'b11, 2'b00, 2'b11, 2'b01, 2'b01, 2'b01, 2'b00, 2'b00, 2'b00, 2'b00, 2'b11, 2'b01, 2'b00, 2'b11, 2'b11, 2'b00, 2'b01, 2'b00, 2'b00, 2'b01, 2'b11, 2'b11, 2'b00, 2'b00, 2'b01, 2'b11, 2'b01, 2'b00, 2'b01 },
		'{ 2'b01, 2'b01, 2'b00, 2'b10, 2'b11, 2'b10, 2'b01, 2'b01, 2'b11, 2'b01, 2'b01, 2'b01, 2'b01, 2'b00, 2'b01, 2'b10, 2'b00, 2'b00, 2'b01, 2'b01, 2'b00, 2'b11, 2'b01, 2'b00, 2'b00, 2'b01, 2'b00, 2'b11, 2'b11, 2'b10, 2'b01, 2'b01, 2'b01, 2'b00, 2'b11, 2'b11, 2'b01, 2'b00, 2'b00, 2'b01, 2'b10, 2'b01, 2'b01, 2'b00, 2'b00, 2'b10, 2'b10, 2'b00, 2'b00, 2'b11, 2'b10, 2'b00, 2'b01, 2'b01, 2'b01, 2'b00, 2'b01, 2'b00, 2'b10, 2'b01, 2'b10, 2'b11, 2'b01, 2'b11 },
		'{ 2'b01, 2'b01, 2'b00, 2'b01, 2'b01, 2'b00, 2'b01, 2'b10, 2'b00, 2'b01, 2'b01, 2'b00, 2'b00, 2'b00, 2'b00, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b00, 2'b01, 2'b00, 2'b11, 2'b00, 2'b00, 2'b01, 2'b11, 2'b01, 2'b01, 2'b01, 2'b00, 2'b11, 2'b01, 2'b11, 2'b01, 2'b01, 2'b10, 2'b00, 2'b10, 2'b00, 2'b01, 2'b00, 2'b11, 2'b11, 2'b00, 2'b11, 2'b00, 2'b11, 2'b00, 2'b10, 2'b10, 2'b11, 2'b10, 2'b01, 2'b00, 2'b00, 2'b01, 2'b00, 2'b00, 2'b00, 2'b10, 2'b10 },
		'{ 2'b00, 2'b00, 2'b01, 2'b01, 2'b01, 2'b00, 2'b01, 2'b11, 2'b00, 2'b01, 2'b10, 2'b00, 2'b00, 2'b10, 2'b00, 2'b01, 2'b11, 2'b00, 2'b01, 2'b00, 2'b01, 2'b01, 2'b00, 2'b11, 2'b00, 2'b11, 2'b00, 2'b11, 2'b00, 2'b01, 2'b10, 2'b00, 2'b01, 2'b01, 2'b11, 2'b01, 2'b10, 2'b01, 2'b00, 2'b01, 2'b01, 2'b11, 2'b01, 2'b00, 2'b01, 2'b01, 2'b11, 2'b01, 2'b11, 2'b01, 2'b00, 2'b00, 2'b00, 2'b00, 2'b11, 2'b01, 2'b00, 2'b01, 2'b00, 2'b11, 2'b01, 2'b10, 2'b01, 2'b00 },
		'{ 2'b00, 2'b00, 2'b11, 2'b00, 2'b01, 2'b01, 2'b00, 2'b01, 2'b00, 2'b00, 2'b11, 2'b01, 2'b00, 2'b11, 2'b01, 2'b10, 2'b00, 2'b00, 2'b00, 2'b01, 2'b01, 2'b11, 2'b11, 2'b11, 2'b00, 2'b11, 2'b00, 2'b01, 2'b00, 2'b01, 2'b11, 2'b11, 2'b01, 2'b00, 2'b01, 2'b00, 2'b00, 2'b11, 2'b01, 2'b01, 2'b11, 2'b01, 2'b00, 2'b10, 2'b01, 2'b00, 2'b11, 2'b01, 2'b10, 2'b11, 2'b11, 2'b00, 2'b10, 2'b00, 2'b00, 2'b01, 2'b01, 2'b00, 2'b00, 2'b01, 2'b00, 2'b10, 2'b01, 2'b01 },
		'{ 2'b01, 2'b00, 2'b01, 2'b11, 2'b00, 2'b01, 2'b11, 2'b00, 2'b00, 2'b10, 2'b11, 2'b01, 2'b01, 2'b00, 2'b01, 2'b00, 2'b00, 2'b00, 2'b11, 2'b00, 2'b01, 2'b10, 2'b01, 2'b01, 2'b00, 2'b11, 2'b01, 2'b00, 2'b00, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b00, 2'b01, 2'b00, 2'b00, 2'b00, 2'b11, 2'b11, 2'b00, 2'b01, 2'b00, 2'b11, 2'b11, 2'b10, 2'b01, 2'b00, 2'b00, 2'b01, 2'b00, 2'b11, 2'b01, 2'b11, 2'b11, 2'b10, 2'b11, 2'b01, 2'b00, 2'b01, 2'b11, 2'b00, 2'b01 },
		'{ 2'b11, 2'b01, 2'b11, 2'b11, 2'b11, 2'b00, 2'b11, 2'b00, 2'b10, 2'b01, 2'b00, 2'b01, 2'b11, 2'b00, 2'b00, 2'b01, 2'b00, 2'b00, 2'b00, 2'b11, 2'b00, 2'b11, 2'b01, 2'b11, 2'b01, 2'b01, 2'b01, 2'b01, 2'b11, 2'b01, 2'b11, 2'b11, 2'b11, 2'b01, 2'b11, 2'b01, 2'b01, 2'b00, 2'b01, 2'b11, 2'b01, 2'b11, 2'b01, 2'b11, 2'b00, 2'b00, 2'b10, 2'b00, 2'b11, 2'b00, 2'b01, 2'b00, 2'b00, 2'b00, 2'b00, 2'b00, 2'b11, 2'b00, 2'b11, 2'b00, 2'b11, 2'b01, 2'b11, 2'b11 },
		'{ 2'b01, 2'b00, 2'b00, 2'b10, 2'b01, 2'b01, 2'b01, 2'b00, 2'b00, 2'b01, 2'b11, 2'b11, 2'b00, 2'b00, 2'b10, 2'b01, 2'b11, 2'b01, 2'b11, 2'b00, 2'b00, 2'b00, 2'b00, 2'b00, 2'b01, 2'b00, 2'b00, 2'b00, 2'b00, 2'b00, 2'b00, 2'b00, 2'b10, 2'b00, 2'b11, 2'b00, 2'b01, 2'b00, 2'b00, 2'b11, 2'b01, 2'b11, 2'b11, 2'b00, 2'b00, 2'b01, 2'b11, 2'b01, 2'b11, 2'b11, 2'b11, 2'b00, 2'b01, 2'b11, 2'b00, 2'b11, 2'b10, 2'b00, 2'b10, 2'b00, 2'b01, 2'b00, 2'b00, 2'b11 },
		'{ 2'b00, 2'b11, 2'b00, 2'b10, 2'b01, 2'b01, 2'b00, 2'b01, 2'b01, 2'b10, 2'b00, 2'b11, 2'b00, 2'b00, 2'b01, 2'b10, 2'b01, 2'b00, 2'b00, 2'b00, 2'b01, 2'b00, 2'b00, 2'b11, 2'b01, 2'b01, 2'b10, 2'b11, 2'b00, 2'b00, 2'b00, 2'b00, 2'b00, 2'b00, 2'b11, 2'b11, 2'b01, 2'b11, 2'b01, 2'b01, 2'b00, 2'b01, 2'b11, 2'b01, 2'b00, 2'b11, 2'b01, 2'b11, 2'b10, 2'b00, 2'b01, 2'b11, 2'b11, 2'b01, 2'b11, 2'b11, 2'b01, 2'b11, 2'b00, 2'b11, 2'b00, 2'b01, 2'b00, 2'b00 },
		'{ 2'b00, 2'b00, 2'b01, 2'b00, 2'b11, 2'b10, 2'b11, 2'b01, 2'b00, 2'b11, 2'b10, 2'b00, 2'b00, 2'b11, 2'b00, 2'b11, 2'b00, 2'b11, 2'b00, 2'b00, 2'b00, 2'b00, 2'b00, 2'b11, 2'b01, 2'b11, 2'b01, 2'b00, 2'b00, 2'b00, 2'b00, 2'b00, 2'b11, 2'b11, 2'b11, 2'b00, 2'b00, 2'b01, 2'b01, 2'b01, 2'b11, 2'b01, 2'b11, 2'b10, 2'b00, 2'b00, 2'b00, 2'b01, 2'b01, 2'b11, 2'b11, 2'b01, 2'b00, 2'b01, 2'b11, 2'b01, 2'b00, 2'b00, 2'b11, 2'b01, 2'b11, 2'b11, 2'b11, 2'b00 },
		'{ 2'b01, 2'b01, 2'b00, 2'b01, 2'b11, 2'b11, 2'b11, 2'b01, 2'b01, 2'b01, 2'b00, 2'b11, 2'b01, 2'b00, 2'b00, 2'b11, 2'b00, 2'b01, 2'b00, 2'b00, 2'b00, 2'b00, 2'b00, 2'b11, 2'b00, 2'b01, 2'b00, 2'b01, 2'b11, 2'b01, 2'b01, 2'b01, 2'b10, 2'b01, 2'b10, 2'b00, 2'b00, 2'b11, 2'b00, 2'b11, 2'b11, 2'b00, 2'b00, 2'b01, 2'b00, 2'b00, 2'b00, 2'b01, 2'b01, 2'b00, 2'b00, 2'b10, 2'b01, 2'b01, 2'b00, 2'b11, 2'b00, 2'b11, 2'b00, 2'b10, 2'b11, 2'b01, 2'b11, 2'b00 },
		'{ 2'b00, 2'b00, 2'b00, 2'b00, 2'b11, 2'b00, 2'b01, 2'b00, 2'b10, 2'b00, 2'b01, 2'b11, 2'b00, 2'b00, 2'b00, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b00, 2'b01, 2'b11, 2'b00, 2'b01, 2'b11, 2'b10, 2'b00, 2'b11, 2'b00, 2'b01, 2'b01, 2'b00, 2'b00, 2'b00, 2'b00, 2'b00, 2'b11, 2'b00, 2'b00, 2'b01, 2'b11, 2'b11, 2'b11, 2'b00, 2'b00, 2'b00, 2'b00, 2'b11, 2'b00, 2'b01, 2'b10, 2'b11, 2'b00, 2'b01, 2'b11, 2'b01, 2'b00, 2'b00, 2'b10, 2'b10, 2'b10, 2'b01, 2'b01 },
		'{ 2'b01, 2'b11, 2'b11, 2'b00, 2'b11, 2'b01, 2'b01, 2'b10, 2'b00, 2'b11, 2'b01, 2'b00, 2'b00, 2'b01, 2'b11, 2'b01, 2'b01, 2'b11, 2'b11, 2'b00, 2'b00, 2'b11, 2'b00, 2'b01, 2'b00, 2'b01, 2'b00, 2'b10, 2'b01, 2'b01, 2'b01, 2'b01, 2'b11, 2'b00, 2'b00, 2'b01, 2'b10, 2'b01, 2'b01, 2'b11, 2'b10, 2'b10, 2'b00, 2'b11, 2'b01, 2'b01, 2'b00, 2'b01, 2'b00, 2'b00, 2'b00, 2'b00, 2'b00, 2'b11, 2'b11, 2'b01, 2'b11, 2'b11, 2'b01, 2'b01, 2'b11, 2'b01, 2'b00, 2'b11 },
		'{ 2'b01, 2'b01, 2'b10, 2'b01, 2'b01, 2'b01, 2'b11, 2'b01, 2'b00, 2'b11, 2'b11, 2'b00, 2'b10, 2'b01, 2'b11, 2'b00, 2'b11, 2'b00, 2'b00, 2'b00, 2'b00, 2'b10, 2'b01, 2'b01, 2'b01, 2'b10, 2'b01, 2'b11, 2'b00, 2'b11, 2'b00, 2'b11, 2'b00, 2'b00, 2'b11, 2'b00, 2'b11, 2'b01, 2'b00, 2'b11, 2'b11, 2'b11, 2'b01, 2'b11, 2'b00, 2'b00, 2'b01, 2'b01, 2'b01, 2'b10, 2'b00, 2'b11, 2'b00, 2'b10, 2'b11, 2'b01, 2'b00, 2'b01, 2'b10, 2'b11, 2'b11, 2'b01, 2'b11, 2'b00 },
		'{ 2'b00, 2'b00, 2'b11, 2'b00, 2'b00, 2'b01, 2'b10, 2'b01, 2'b00, 2'b01, 2'b10, 2'b00, 2'b01, 2'b11, 2'b11, 2'b00, 2'b11, 2'b00, 2'b01, 2'b10, 2'b00, 2'b10, 2'b11, 2'b00, 2'b10, 2'b11, 2'b01, 2'b11, 2'b00, 2'b01, 2'b00, 2'b11, 2'b01, 2'b00, 2'b00, 2'b00, 2'b01, 2'b01, 2'b10, 2'b00, 2'b01, 2'b00, 2'b00, 2'b11, 2'b00, 2'b00, 2'b01, 2'b00, 2'b01, 2'b01, 2'b01, 2'b00, 2'b01, 2'b00, 2'b11, 2'b10, 2'b00, 2'b11, 2'b01, 2'b11, 2'b01, 2'b01, 2'b01, 2'b01 },
		'{ 2'b01, 2'b10, 2'b01, 2'b00, 2'b00, 2'b01, 2'b11, 2'b01, 2'b11, 2'b10, 2'b11, 2'b00, 2'b00, 2'b00, 2'b00, 2'b00, 2'b01, 2'b10, 2'b11, 2'b11, 2'b01, 2'b01, 2'b01, 2'b11, 2'b00, 2'b01, 2'b01, 2'b00, 2'b11, 2'b00, 2'b00, 2'b11, 2'b01, 2'b00, 2'b11, 2'b00, 2'b01, 2'b11, 2'b01, 2'b01, 2'b01, 2'b11, 2'b11, 2'b00, 2'b11, 2'b01, 2'b00, 2'b11, 2'b11, 2'b01, 2'b00, 2'b01, 2'b00, 2'b11, 2'b11, 2'b11, 2'b01, 2'b00, 2'b00, 2'b00, 2'b00, 2'b11, 2'b01, 2'b01 },
		'{ 2'b00, 2'b01, 2'b01, 2'b01, 2'b11, 2'b01, 2'b01, 2'b10, 2'b11, 2'b00, 2'b11, 2'b00, 2'b00, 2'b11, 2'b00, 2'b00, 2'b00, 2'b11, 2'b01, 2'b01, 2'b01, 2'b00, 2'b11, 2'b00, 2'b01, 2'b00, 2'b00, 2'b11, 2'b00, 2'b00, 2'b10, 2'b00, 2'b00, 2'b00, 2'b00, 2'b00, 2'b11, 2'b11, 2'b11, 2'b11, 2'b11, 2'b01, 2'b01, 2'b11, 2'b11, 2'b00, 2'b11, 2'b11, 2'b00, 2'b01, 2'b01, 2'b01, 2'b10, 2'b00, 2'b01, 2'b00, 2'b11, 2'b01, 2'b00, 2'b01, 2'b11, 2'b01, 2'b00, 2'b00 },
		'{ 2'b01, 2'b00, 2'b11, 2'b11, 2'b10, 2'b01, 2'b11, 2'b00, 2'b01, 2'b01, 2'b00, 2'b01, 2'b01, 2'b11, 2'b00, 2'b00, 2'b00, 2'b11, 2'b00, 2'b11, 2'b11, 2'b00, 2'b00, 2'b00, 2'b01, 2'b00, 2'b01, 2'b00, 2'b00, 2'b11, 2'b00, 2'b01, 2'b11, 2'b00, 2'b11, 2'b00, 2'b11, 2'b00, 2'b01, 2'b00, 2'b10, 2'b11, 2'b01, 2'b11, 2'b00, 2'b00, 2'b11, 2'b11, 2'b00, 2'b00, 2'b00, 2'b01, 2'b11, 2'b00, 2'b10, 2'b01, 2'b01, 2'b11, 2'b00, 2'b11, 2'b00, 2'b11, 2'b01, 2'b00 },
		'{ 2'b10, 2'b00, 2'b00, 2'b00, 2'b01, 2'b00, 2'b01, 2'b10, 2'b00, 2'b11, 2'b01, 2'b00, 2'b00, 2'b11, 2'b11, 2'b00, 2'b11, 2'b00, 2'b10, 2'b01, 2'b01, 2'b11, 2'b01, 2'b11, 2'b00, 2'b11, 2'b00, 2'b00, 2'b11, 2'b01, 2'b11, 2'b00, 2'b00, 2'b00, 2'b00, 2'b01, 2'b00, 2'b10, 2'b00, 2'b11, 2'b01, 2'b00, 2'b00, 2'b01, 2'b10, 2'b01, 2'b01, 2'b11, 2'b01, 2'b00, 2'b00, 2'b11, 2'b00, 2'b11, 2'b00, 2'b10, 2'b01, 2'b00, 2'b11, 2'b01, 2'b10, 2'b00, 2'b00, 2'b01 },
		'{ 2'b00, 2'b11, 2'b00, 2'b11, 2'b11, 2'b01, 2'b00, 2'b11, 2'b01, 2'b11, 2'b00, 2'b11, 2'b01, 2'b00, 2'b01, 2'b01, 2'b00, 2'b01, 2'b00, 2'b00, 2'b11, 2'b01, 2'b00, 2'b11, 2'b11, 2'b00, 2'b00, 2'b00, 2'b01, 2'b00, 2'b00, 2'b00, 2'b01, 2'b00, 2'b11, 2'b00, 2'b00, 2'b11, 2'b01, 2'b01, 2'b00, 2'b11, 2'b01, 2'b11, 2'b11, 2'b01, 2'b00, 2'b11, 2'b00, 2'b01, 2'b00, 2'b00, 2'b01, 2'b10, 2'b01, 2'b00, 2'b01, 2'b01, 2'b01, 2'b11, 2'b01, 2'b00, 2'b01, 2'b01 },
		'{ 2'b01, 2'b00, 2'b01, 2'b11, 2'b00, 2'b10, 2'b11, 2'b11, 2'b00, 2'b01, 2'b00, 2'b10, 2'b01, 2'b11, 2'b11, 2'b00, 2'b11, 2'b00, 2'b11, 2'b11, 2'b00, 2'b01, 2'b00, 2'b00, 2'b01, 2'b11, 2'b01, 2'b11, 2'b00, 2'b00, 2'b01, 2'b11, 2'b11, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b00, 2'b00, 2'b00, 2'b01, 2'b01, 2'b00, 2'b01, 2'b11, 2'b01, 2'b01, 2'b00, 2'b00, 2'b01, 2'b11, 2'b11, 2'b00, 2'b11, 2'b00, 2'b01, 2'b11, 2'b01, 2'b01, 2'b11, 2'b00, 2'b01, 2'b10 },
		'{ 2'b01, 2'b00, 2'b11, 2'b00, 2'b00, 2'b00, 2'b11, 2'b00, 2'b00, 2'b00, 2'b00, 2'b11, 2'b00, 2'b00, 2'b01, 2'b11, 2'b10, 2'b11, 2'b01, 2'b01, 2'b11, 2'b00, 2'b01, 2'b00, 2'b00, 2'b01, 2'b00, 2'b00, 2'b00, 2'b01, 2'b00, 2'b01, 2'b01, 2'b00, 2'b01, 2'b11, 2'b11, 2'b11, 2'b00, 2'b01, 2'b01, 2'b01, 2'b11, 2'b11, 2'b01, 2'b00, 2'b11, 2'b00, 2'b00, 2'b10, 2'b11, 2'b11, 2'b01, 2'b01, 2'b01, 2'b10, 2'b01, 2'b00, 2'b01, 2'b10, 2'b11, 2'b11, 2'b01, 2'b01 },
		'{ 2'b11, 2'b11, 2'b10, 2'b01, 2'b11, 2'b01, 2'b11, 2'b01, 2'b11, 2'b01, 2'b01, 2'b11, 2'b01, 2'b01, 2'b00, 2'b00, 2'b01, 2'b00, 2'b00, 2'b11, 2'b11, 2'b11, 2'b01, 2'b10, 2'b00, 2'b01, 2'b00, 2'b00, 2'b00, 2'b00, 2'b11, 2'b00, 2'b11, 2'b10, 2'b01, 2'b11, 2'b01, 2'b10, 2'b01, 2'b00, 2'b00, 2'b11, 2'b01, 2'b10, 2'b01, 2'b00, 2'b01, 2'b00, 2'b01, 2'b01, 2'b00, 2'b00, 2'b00, 2'b11, 2'b11, 2'b11, 2'b11, 2'b11, 2'b11, 2'b01, 2'b10, 2'b11, 2'b11, 2'b00 },
		'{ 2'b11, 2'b11, 2'b00, 2'b00, 2'b00, 2'b01, 2'b01, 2'b00, 2'b01, 2'b01, 2'b11, 2'b01, 2'b00, 2'b01, 2'b01, 2'b01, 2'b10, 2'b11, 2'b11, 2'b01, 2'b00, 2'b00, 2'b11, 2'b00, 2'b00, 2'b11, 2'b11, 2'b00, 2'b00, 2'b00, 2'b00, 2'b10, 2'b00, 2'b00, 2'b00, 2'b10, 2'b00, 2'b10, 2'b00, 2'b01, 2'b01, 2'b00, 2'b00, 2'b00, 2'b01, 2'b00, 2'b00, 2'b00, 2'b11, 2'b00, 2'b01, 2'b00, 2'b01, 2'b11, 2'b01, 2'b00, 2'b01, 2'b00, 2'b11, 2'b00, 2'b11, 2'b11, 2'b11, 2'b00 }
	};
    
endpackage