//===========================================================
// Purpose: Segmentation package
// Used in: image_segmentation
//===========================================================
package segmentation_pkg;
  typedef enum bit {IDLE, TRANSMIT} states_t;
endpackage