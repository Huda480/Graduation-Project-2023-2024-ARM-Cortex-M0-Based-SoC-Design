library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
library UNISIM;
use UNISIM.VCOMPONENTS.ALL;
use UNISIM.VPKG.ALL;

entity FFT is
  port (
    clk : in STD_LOGIC := 'X'; 
    ce : in STD_LOGIC := 'X'; 
    start : in STD_LOGIC := 'X'; 
    cp_len_we : in STD_LOGIC := 'X'; 
    fwd_inv : in STD_LOGIC := 'X'; 
    fwd_inv_we : in STD_LOGIC := 'X'; 
    scale_sch_we : in STD_LOGIC := 'X'; 
    rfd : out STD_LOGIC; 
    busy : out STD_LOGIC; 
    edone : out STD_LOGIC; 
    done : out STD_LOGIC; 
    dv : out STD_LOGIC; 
    cpv : out STD_LOGIC; 
    rfs : out STD_LOGIC; 
    cp_len : in STD_LOGIC_VECTOR ( 5 downto 0 ); 
    xn_re : in STD_LOGIC_VECTOR ( 11 downto 0 ); 
    xn_im : in STD_LOGIC_VECTOR ( 11 downto 0 ); 
    scale_sch : in STD_LOGIC_VECTOR ( 5 downto 0 ); 
    xn_index : out STD_LOGIC_VECTOR ( 5 downto 0 ); 
    xk_index : out STD_LOGIC_VECTOR ( 5 downto 0 ); 
    xk_re : out STD_LOGIC_VECTOR ( 11 downto 0 ); 
    xk_im : out STD_LOGIC_VECTOR ( 11 downto 0 ) 
  );
  attribute dont_touch : string;
attribute dont_touch of FFT : entity is "true|yes";
end FFT;
architecture STRUCTURE of FFT is
--attribute dont_touch : string;
attribute dont_touch of STRUCTURE : architecture is "yes";
  signal NlwRenamedSig_OI_U0_i_synth_non_floating_point_arch_d_xfft_inst_FLOW_load_enable : STD_LOGIC; 
  signal U0_i_synth_non_floating_point_arch_d_xfft_inst_has_bit_reverse_busy_gen_busy_i : STD_LOGIC; 
  signal NlwRenamedSig_OI_U0_i_synth_non_floating_point_arch_d_xfft_inst_done_int_d : STD_LOGIC; 
  signal U0_i_synth_non_floating_point_arch_d_xfft_inst_DONE : STD_LOGIC; 
  signal U0_i_synth_non_floating_point_arch_d_xfft_inst_DV : STD_LOGIC; 
  signal NlwRenamedSig_OI_cpv : STD_LOGIC; 
  signal NlwRenamedSig_OI_rfs : STD_LOGIC; 
  signal sig00000001 : STD_LOGIC; 
  signal sig00000002 : STD_LOGIC; 
  signal sig00000003 : STD_LOGIC; 
  signal sig00000004 : STD_LOGIC; 
  signal sig00000005 : STD_LOGIC; 
  signal sig00000006 : STD_LOGIC; 
  signal sig00000007 : STD_LOGIC; 
  signal sig00000008 : STD_LOGIC; 
  signal sig00000009 : STD_LOGIC; 
  signal sig0000000a : STD_LOGIC; 
  signal sig0000000b : STD_LOGIC; 
  signal sig0000000c : STD_LOGIC; 
  signal sig0000000d : STD_LOGIC; 
  signal sig0000000e : STD_LOGIC; 
  signal sig0000000f : STD_LOGIC; 
  signal sig00000010 : STD_LOGIC; 
  signal sig00000011 : STD_LOGIC; 
  signal sig00000012 : STD_LOGIC; 
  signal sig00000013 : STD_LOGIC; 
  signal sig00000014 : STD_LOGIC; 
  signal sig00000015 : STD_LOGIC; 
  signal sig00000016 : STD_LOGIC; 
  signal sig00000017 : STD_LOGIC; 
  signal sig00000018 : STD_LOGIC; 
  signal sig00000019 : STD_LOGIC; 
  signal sig0000001a : STD_LOGIC; 
  signal sig0000001b : STD_LOGIC; 
  signal sig0000001c : STD_LOGIC; 
  signal sig0000001d : STD_LOGIC; 
  signal sig0000001e : STD_LOGIC; 
  signal sig0000001f : STD_LOGIC; 
  signal sig00000020 : STD_LOGIC; 
  signal sig00000021 : STD_LOGIC; 
  signal sig00000022 : STD_LOGIC; 
  signal sig00000023 : STD_LOGIC; 
  signal sig00000024 : STD_LOGIC; 
  signal sig00000025 : STD_LOGIC; 
  signal sig00000026 : STD_LOGIC; 
  signal sig00000027 : STD_LOGIC; 
  signal sig00000028 : STD_LOGIC; 
  signal sig00000029 : STD_LOGIC; 
  signal sig0000002a : STD_LOGIC; 
  signal sig0000002b : STD_LOGIC; 
  signal sig0000002c : STD_LOGIC; 
  signal sig0000002d : STD_LOGIC; 
  signal sig0000002e : STD_LOGIC; 
  signal sig0000002f : STD_LOGIC; 
  signal sig00000030 : STD_LOGIC; 
  signal sig00000031 : STD_LOGIC; 
  signal sig00000032 : STD_LOGIC; 
  signal sig00000033 : STD_LOGIC; 
  signal sig00000034 : STD_LOGIC; 
  signal sig00000035 : STD_LOGIC; 
  signal sig00000036 : STD_LOGIC; 
  signal sig00000037 : STD_LOGIC; 
  signal sig00000038 : STD_LOGIC; 
  signal sig00000039 : STD_LOGIC; 
  signal sig0000003a : STD_LOGIC; 
  signal sig0000003b : STD_LOGIC; 
  signal sig0000003c : STD_LOGIC; 
  signal sig0000003d : STD_LOGIC; 
  signal sig0000003e : STD_LOGIC; 
  signal sig0000003f : STD_LOGIC; 
  signal sig00000040 : STD_LOGIC; 
  signal sig00000041 : STD_LOGIC; 
  signal sig00000042 : STD_LOGIC; 
  signal sig00000043 : STD_LOGIC; 
  signal sig00000044 : STD_LOGIC; 
  signal sig00000045 : STD_LOGIC; 
  signal sig00000046 : STD_LOGIC; 
  signal sig00000047 : STD_LOGIC; 
  signal sig00000048 : STD_LOGIC; 
  signal sig00000049 : STD_LOGIC; 
  signal sig0000004a : STD_LOGIC; 
  signal sig0000004b : STD_LOGIC; 
  signal sig0000004c : STD_LOGIC; 
  signal sig0000004d : STD_LOGIC; 
  signal sig0000004e : STD_LOGIC; 
  signal sig0000004f : STD_LOGIC; 
  signal sig00000050 : STD_LOGIC; 
  signal sig00000051 : STD_LOGIC; 
  signal sig00000052 : STD_LOGIC; 
  signal sig00000053 : STD_LOGIC; 
  signal sig00000054 : STD_LOGIC; 
  signal sig00000055 : STD_LOGIC; 
  signal sig00000056 : STD_LOGIC; 
  signal sig00000057 : STD_LOGIC; 
  signal sig00000058 : STD_LOGIC; 
  signal sig00000059 : STD_LOGIC; 
  signal sig0000005a : STD_LOGIC; 
  signal sig0000005b : STD_LOGIC; 
  signal sig0000005c : STD_LOGIC; 
  signal sig0000005d : STD_LOGIC; 
  signal sig0000005e : STD_LOGIC; 
  signal sig0000005f : STD_LOGIC; 
  signal sig00000060 : STD_LOGIC; 
  signal sig00000061 : STD_LOGIC; 
  signal sig00000062 : STD_LOGIC; 
  signal sig00000063 : STD_LOGIC; 
  signal sig00000064 : STD_LOGIC; 
  signal sig00000065 : STD_LOGIC; 
  signal sig00000066 : STD_LOGIC; 
  signal sig00000067 : STD_LOGIC; 
  signal sig00000068 : STD_LOGIC; 
  signal sig00000069 : STD_LOGIC; 
  signal sig0000006a : STD_LOGIC; 
  signal sig0000006b : STD_LOGIC; 
  signal sig0000006c : STD_LOGIC; 
  signal sig0000006d : STD_LOGIC; 
  signal sig0000006e : STD_LOGIC; 
  signal sig0000006f : STD_LOGIC; 
  signal sig00000070 : STD_LOGIC; 
  signal sig00000071 : STD_LOGIC; 
  signal sig00000072 : STD_LOGIC; 
  signal sig00000073 : STD_LOGIC; 
  signal sig00000074 : STD_LOGIC; 
  signal sig00000075 : STD_LOGIC; 
  signal sig00000076 : STD_LOGIC; 
  signal sig00000077 : STD_LOGIC; 
  signal sig00000078 : STD_LOGIC; 
  signal sig00000079 : STD_LOGIC; 
  signal sig0000007a : STD_LOGIC; 
  signal sig0000007b : STD_LOGIC; 
  signal sig0000007c : STD_LOGIC; 
  signal sig0000007d : STD_LOGIC; 
  signal sig0000007e : STD_LOGIC; 
  signal sig0000007f : STD_LOGIC; 
  signal sig00000080 : STD_LOGIC; 
  signal sig00000081 : STD_LOGIC; 
  signal sig00000082 : STD_LOGIC; 
  signal sig00000083 : STD_LOGIC; 
  signal sig00000084 : STD_LOGIC; 
  signal sig00000085 : STD_LOGIC; 
  signal sig00000086 : STD_LOGIC; 
  signal sig00000087 : STD_LOGIC; 
  signal sig00000088 : STD_LOGIC; 
  signal sig00000089 : STD_LOGIC; 
  signal sig0000008a : STD_LOGIC; 
  signal sig0000008b : STD_LOGIC; 
  signal sig0000008c : STD_LOGIC; 
  signal sig0000008d : STD_LOGIC; 
  signal sig0000008e : STD_LOGIC; 
  signal sig0000008f : STD_LOGIC; 
  signal sig00000090 : STD_LOGIC; 
  signal sig00000091 : STD_LOGIC; 
  signal sig00000092 : STD_LOGIC; 
  signal sig00000093 : STD_LOGIC; 
  signal sig00000094 : STD_LOGIC; 
  signal sig00000095 : STD_LOGIC; 
  signal sig00000096 : STD_LOGIC; 
  signal sig00000097 : STD_LOGIC; 
  signal sig00000098 : STD_LOGIC; 
  signal sig00000099 : STD_LOGIC; 
  signal sig0000009a : STD_LOGIC; 
  signal sig0000009b : STD_LOGIC; 
  signal sig0000009c : STD_LOGIC; 
  signal sig0000009d : STD_LOGIC; 
  signal sig0000009e : STD_LOGIC; 
  signal sig0000009f : STD_LOGIC; 
  signal sig000000a0 : STD_LOGIC; 
  signal sig000000a1 : STD_LOGIC; 
  signal sig000000a2 : STD_LOGIC; 
  signal sig000000a3 : STD_LOGIC; 
  signal sig000000a4 : STD_LOGIC; 
  signal sig000000a5 : STD_LOGIC; 
  signal sig000000a6 : STD_LOGIC; 
  signal sig000000a7 : STD_LOGIC; 
  signal sig000000a8 : STD_LOGIC; 
  signal sig000000a9 : STD_LOGIC; 
  signal sig000000aa : STD_LOGIC; 
  signal sig000000ab : STD_LOGIC; 
  signal sig000000ac : STD_LOGIC; 
  signal sig000000ad : STD_LOGIC; 
  signal sig000000ae : STD_LOGIC; 
  signal sig000000af : STD_LOGIC; 
  signal sig000000b0 : STD_LOGIC; 
  signal sig000000b1 : STD_LOGIC; 
  signal sig000000b2 : STD_LOGIC; 
  signal sig000000b3 : STD_LOGIC; 
  signal sig000000b4 : STD_LOGIC; 
  signal sig000000b5 : STD_LOGIC; 
  signal sig000000b6 : STD_LOGIC; 
  signal sig000000b7 : STD_LOGIC; 
  signal sig000000b8 : STD_LOGIC; 
  signal sig000000b9 : STD_LOGIC; 
  signal sig000000ba : STD_LOGIC; 
  signal sig000000bb : STD_LOGIC; 
  signal sig000000bc : STD_LOGIC; 
  signal sig000000bd : STD_LOGIC; 
  signal sig000000be : STD_LOGIC; 
  signal sig000000bf : STD_LOGIC; 
  signal sig000000c0 : STD_LOGIC; 
  signal sig000000c1 : STD_LOGIC; 
  signal sig000000c2 : STD_LOGIC; 
  signal sig000000c3 : STD_LOGIC; 
  signal sig000000c4 : STD_LOGIC; 
  signal sig000000c5 : STD_LOGIC; 
  signal sig000000c6 : STD_LOGIC; 
  signal sig000000c7 : STD_LOGIC; 
  signal sig000000c8 : STD_LOGIC; 
  signal sig000000c9 : STD_LOGIC; 
  signal sig000000ca : STD_LOGIC; 
  signal sig000000cb : STD_LOGIC; 
  signal sig000000cc : STD_LOGIC; 
  signal sig000000cd : STD_LOGIC; 
  signal sig000000ce : STD_LOGIC; 
  signal sig000000cf : STD_LOGIC; 
  signal sig000000d0 : STD_LOGIC; 
  signal sig000000d1 : STD_LOGIC; 
  signal sig000000d2 : STD_LOGIC; 
  signal sig000000d3 : STD_LOGIC; 
  signal sig000000d4 : STD_LOGIC; 
  signal sig000000d5 : STD_LOGIC; 
  signal sig000000d6 : STD_LOGIC; 
  signal sig000000d7 : STD_LOGIC; 
  signal sig000000d8 : STD_LOGIC; 
  signal sig000000d9 : STD_LOGIC; 
  signal sig000000da : STD_LOGIC; 
  signal sig000000db : STD_LOGIC; 
  signal sig000000dc : STD_LOGIC; 
  signal sig000000dd : STD_LOGIC; 
  signal sig000000de : STD_LOGIC; 
  signal sig000000df : STD_LOGIC; 
  signal sig000000e0 : STD_LOGIC; 
  signal sig000000e1 : STD_LOGIC; 
  signal sig000000e2 : STD_LOGIC; 
  signal sig000000e3 : STD_LOGIC; 
  signal sig000000e4 : STD_LOGIC; 
  signal sig000000e5 : STD_LOGIC; 
  signal sig000000e6 : STD_LOGIC; 
  signal sig000000e7 : STD_LOGIC; 
  signal sig000000e8 : STD_LOGIC; 
  signal sig000000e9 : STD_LOGIC; 
  signal sig000000ea : STD_LOGIC; 
  signal sig000000eb : STD_LOGIC; 
  signal sig000000ec : STD_LOGIC; 
  signal sig000000ed : STD_LOGIC; 
  signal sig000000ee : STD_LOGIC; 
  signal sig000000ef : STD_LOGIC; 
  signal sig000000f0 : STD_LOGIC; 
  signal sig000000f1 : STD_LOGIC; 
  signal sig000000f2 : STD_LOGIC; 
  signal sig000000f3 : STD_LOGIC; 
  signal sig000000f4 : STD_LOGIC; 
  signal sig000000f5 : STD_LOGIC; 
  signal sig000000f6 : STD_LOGIC; 
  signal sig000000f7 : STD_LOGIC; 
  signal sig000000f8 : STD_LOGIC; 
  signal sig000000f9 : STD_LOGIC; 
  signal sig000000fa : STD_LOGIC; 
  signal sig000000fb : STD_LOGIC; 
  signal sig000000fc : STD_LOGIC; 
  signal sig000000fd : STD_LOGIC; 
  signal sig000000fe : STD_LOGIC; 
  signal sig000000ff : STD_LOGIC; 
  signal sig00000100 : STD_LOGIC; 
  signal sig00000101 : STD_LOGIC; 
  signal sig00000102 : STD_LOGIC; 
  signal sig00000103 : STD_LOGIC; 
  signal sig00000104 : STD_LOGIC; 
  signal sig00000105 : STD_LOGIC; 
  signal sig00000106 : STD_LOGIC; 
  signal sig00000107 : STD_LOGIC; 
  signal sig00000108 : STD_LOGIC; 
  signal sig00000109 : STD_LOGIC; 
  signal sig0000010a : STD_LOGIC; 
  signal sig0000010b : STD_LOGIC; 
  signal sig0000010c : STD_LOGIC; 
  signal sig0000010d : STD_LOGIC; 
  signal sig0000010e : STD_LOGIC; 
  signal sig0000010f : STD_LOGIC; 
  signal sig00000110 : STD_LOGIC; 
  signal sig00000111 : STD_LOGIC; 
  signal sig00000112 : STD_LOGIC; 
  signal sig00000113 : STD_LOGIC; 
  signal sig00000114 : STD_LOGIC; 
  signal sig00000115 : STD_LOGIC; 
  signal sig00000116 : STD_LOGIC; 
  signal sig00000117 : STD_LOGIC; 
  signal sig00000118 : STD_LOGIC; 
  signal sig00000119 : STD_LOGIC; 
  signal sig0000011a : STD_LOGIC; 
  signal sig0000011b : STD_LOGIC; 
  signal sig0000011c : STD_LOGIC; 
  signal sig0000011d : STD_LOGIC; 
  signal sig0000011e : STD_LOGIC; 
  signal sig0000011f : STD_LOGIC; 
  signal sig00000120 : STD_LOGIC; 
  signal sig00000121 : STD_LOGIC; 
  signal sig00000122 : STD_LOGIC; 
  signal sig00000123 : STD_LOGIC; 
  signal sig00000124 : STD_LOGIC; 
  signal sig00000125 : STD_LOGIC; 
  signal sig00000126 : STD_LOGIC; 
  signal sig00000127 : STD_LOGIC; 
  signal sig00000128 : STD_LOGIC; 
  signal sig00000129 : STD_LOGIC; 
  signal sig0000012a : STD_LOGIC; 
  signal sig0000012b : STD_LOGIC; 
  signal sig0000012c : STD_LOGIC; 
  signal sig0000012d : STD_LOGIC; 
  signal sig0000012e : STD_LOGIC; 
  signal sig0000012f : STD_LOGIC; 
  signal sig00000130 : STD_LOGIC; 
  signal sig00000131 : STD_LOGIC; 
  signal sig00000132 : STD_LOGIC; 
  signal sig00000133 : STD_LOGIC; 
  signal sig00000134 : STD_LOGIC; 
  signal sig00000135 : STD_LOGIC; 
  signal sig00000136 : STD_LOGIC; 
  signal sig00000137 : STD_LOGIC; 
  signal sig00000138 : STD_LOGIC; 
  signal sig00000139 : STD_LOGIC; 
  signal sig0000013a : STD_LOGIC; 
  signal sig0000013b : STD_LOGIC; 
  signal sig0000013c : STD_LOGIC; 
  signal sig0000013d : STD_LOGIC; 
  signal sig0000013e : STD_LOGIC; 
  signal sig0000013f : STD_LOGIC; 
  signal sig00000140 : STD_LOGIC; 
  signal sig00000141 : STD_LOGIC; 
  signal sig00000142 : STD_LOGIC; 
  signal sig00000143 : STD_LOGIC; 
  signal sig00000144 : STD_LOGIC; 
  signal sig00000145 : STD_LOGIC; 
  signal sig00000146 : STD_LOGIC; 
  signal sig00000147 : STD_LOGIC; 
  signal sig00000148 : STD_LOGIC; 
  signal sig00000149 : STD_LOGIC; 
  signal sig0000014a : STD_LOGIC; 
  signal sig0000014b : STD_LOGIC; 
  signal sig0000014c : STD_LOGIC; 
  signal sig0000014d : STD_LOGIC; 
  signal sig0000014e : STD_LOGIC; 
  signal sig0000014f : STD_LOGIC; 
  signal sig00000150 : STD_LOGIC; 
  signal sig00000151 : STD_LOGIC; 
  signal sig00000152 : STD_LOGIC; 
  signal sig00000153 : STD_LOGIC; 
  signal sig00000154 : STD_LOGIC; 
  signal sig00000155 : STD_LOGIC; 
  signal sig00000156 : STD_LOGIC; 
  signal sig00000157 : STD_LOGIC; 
  signal sig00000158 : STD_LOGIC; 
  signal sig00000159 : STD_LOGIC; 
  signal sig0000015a : STD_LOGIC; 
  signal sig0000015b : STD_LOGIC; 
  signal sig0000015c : STD_LOGIC; 
  signal sig0000015d : STD_LOGIC; 
  signal sig0000015e : STD_LOGIC; 
  signal sig0000015f : STD_LOGIC; 
  signal sig00000160 : STD_LOGIC; 
  signal sig00000161 : STD_LOGIC; 
  signal sig00000162 : STD_LOGIC; 
  signal sig00000163 : STD_LOGIC; 
  signal sig00000164 : STD_LOGIC; 
  signal sig00000165 : STD_LOGIC; 
  signal sig00000166 : STD_LOGIC; 
  signal sig00000167 : STD_LOGIC; 
  signal sig00000168 : STD_LOGIC; 
  signal sig00000169 : STD_LOGIC; 
  signal sig0000016a : STD_LOGIC; 
  signal sig0000016b : STD_LOGIC; 
  signal sig0000016c : STD_LOGIC; 
  signal sig0000016d : STD_LOGIC; 
  signal sig0000016e : STD_LOGIC; 
  signal sig0000016f : STD_LOGIC; 
  signal sig00000170 : STD_LOGIC; 
  signal sig00000171 : STD_LOGIC; 
  signal sig00000172 : STD_LOGIC; 
  signal sig00000173 : STD_LOGIC; 
  signal sig00000174 : STD_LOGIC; 
  signal sig00000175 : STD_LOGIC; 
  signal sig00000176 : STD_LOGIC; 
  signal sig00000177 : STD_LOGIC; 
  signal sig00000178 : STD_LOGIC; 
  signal sig00000179 : STD_LOGIC; 
  signal sig0000017a : STD_LOGIC; 
  signal sig0000017b : STD_LOGIC; 
  signal sig0000017c : STD_LOGIC; 
  signal sig0000017d : STD_LOGIC; 
  signal sig0000017e : STD_LOGIC; 
  signal sig0000017f : STD_LOGIC; 
  signal sig00000180 : STD_LOGIC; 
  signal sig00000181 : STD_LOGIC; 
  signal sig00000182 : STD_LOGIC; 
  signal sig00000183 : STD_LOGIC; 
  signal sig00000184 : STD_LOGIC; 
  signal sig00000185 : STD_LOGIC; 
  signal sig00000186 : STD_LOGIC; 
  signal sig00000187 : STD_LOGIC; 
  signal sig00000188 : STD_LOGIC; 
  signal sig00000189 : STD_LOGIC; 
  signal sig0000018a : STD_LOGIC; 
  signal sig0000018b : STD_LOGIC; 
  signal sig0000018c : STD_LOGIC; 
  signal sig0000018d : STD_LOGIC; 
  signal sig0000018e : STD_LOGIC; 
  signal sig0000018f : STD_LOGIC; 
  signal sig00000190 : STD_LOGIC; 
  signal sig00000191 : STD_LOGIC; 
  signal sig00000192 : STD_LOGIC; 
  signal sig00000193 : STD_LOGIC; 
  signal sig00000194 : STD_LOGIC; 
  signal sig00000195 : STD_LOGIC; 
  signal sig00000196 : STD_LOGIC; 
  signal sig00000197 : STD_LOGIC; 
  signal sig00000198 : STD_LOGIC; 
  signal sig00000199 : STD_LOGIC; 
  signal sig0000019a : STD_LOGIC; 
  signal sig0000019b : STD_LOGIC; 
  signal sig0000019c : STD_LOGIC; 
  signal sig0000019d : STD_LOGIC; 
  signal sig0000019e : STD_LOGIC; 
  signal sig0000019f : STD_LOGIC; 
  signal sig000001a0 : STD_LOGIC; 
  signal sig000001a1 : STD_LOGIC; 
  signal sig000001a2 : STD_LOGIC; 
  signal sig000001a3 : STD_LOGIC; 
  signal sig000001a4 : STD_LOGIC; 
  signal sig000001a5 : STD_LOGIC; 
  signal sig000001a6 : STD_LOGIC; 
  signal sig000001a7 : STD_LOGIC; 
  signal sig000001a8 : STD_LOGIC; 
  signal sig000001a9 : STD_LOGIC; 
  signal sig000001aa : STD_LOGIC; 
  signal sig000001ab : STD_LOGIC; 
  signal sig000001ac : STD_LOGIC; 
  signal sig000001ad : STD_LOGIC; 
  signal sig000001ae : STD_LOGIC; 
  signal sig000001af : STD_LOGIC; 
  signal sig000001b0 : STD_LOGIC; 
  signal sig000001b1 : STD_LOGIC; 
  signal sig000001b2 : STD_LOGIC; 
  signal sig000001b3 : STD_LOGIC; 
  signal sig000001b4 : STD_LOGIC; 
  signal sig000001b5 : STD_LOGIC; 
  signal sig000001b6 : STD_LOGIC; 
  signal sig000001b7 : STD_LOGIC; 
  signal sig000001b8 : STD_LOGIC; 
  signal sig000001b9 : STD_LOGIC; 
  signal sig000001ba : STD_LOGIC; 
  signal sig000001bb : STD_LOGIC; 
  signal sig000001bc : STD_LOGIC; 
  signal sig000001bd : STD_LOGIC; 
  signal sig000001be : STD_LOGIC; 
  signal sig000001bf : STD_LOGIC; 
  signal sig000001c0 : STD_LOGIC; 
  signal sig000001c1 : STD_LOGIC; 
  signal sig000001c2 : STD_LOGIC; 
  signal sig000001c3 : STD_LOGIC; 
  signal sig000001c4 : STD_LOGIC; 
  signal sig000001c5 : STD_LOGIC; 
  signal sig000001c6 : STD_LOGIC; 
  signal sig000001c7 : STD_LOGIC; 
  signal sig000001c8 : STD_LOGIC; 
  signal sig000001c9 : STD_LOGIC; 
  signal sig000001ca : STD_LOGIC; 
  signal sig000001cb : STD_LOGIC; 
  signal sig000001cc : STD_LOGIC; 
  signal sig000001cd : STD_LOGIC; 
  signal sig000001ce : STD_LOGIC; 
  signal sig000001cf : STD_LOGIC; 
  signal sig000001d0 : STD_LOGIC; 
  signal sig000001d1 : STD_LOGIC; 
  signal sig000001d2 : STD_LOGIC; 
  signal sig000001d3 : STD_LOGIC; 
  signal sig000001d4 : STD_LOGIC; 
  signal sig000001d5 : STD_LOGIC; 
  signal sig000001d6 : STD_LOGIC; 
  signal sig000001d7 : STD_LOGIC; 
  signal sig000001d8 : STD_LOGIC; 
  signal sig000001d9 : STD_LOGIC; 
  signal sig000001da : STD_LOGIC; 
  signal sig000001db : STD_LOGIC; 
  signal sig000001dc : STD_LOGIC; 
  signal sig000001dd : STD_LOGIC; 
  signal sig000001de : STD_LOGIC; 
  signal sig000001df : STD_LOGIC; 
  signal sig000001e0 : STD_LOGIC; 
  signal sig000001e1 : STD_LOGIC; 
  signal sig000001e2 : STD_LOGIC; 
  signal sig000001e3 : STD_LOGIC; 
  signal sig000001e4 : STD_LOGIC; 
  signal sig000001e5 : STD_LOGIC; 
  signal sig000001e6 : STD_LOGIC; 
  signal sig000001e7 : STD_LOGIC; 
  signal sig000001e8 : STD_LOGIC; 
  signal sig000001e9 : STD_LOGIC; 
  signal sig000001ea : STD_LOGIC; 
  signal sig000001eb : STD_LOGIC; 
  signal sig000001ec : STD_LOGIC; 
  signal sig000001ed : STD_LOGIC; 
  signal sig000001ee : STD_LOGIC; 
  signal sig000001ef : STD_LOGIC; 
  signal sig000001f0 : STD_LOGIC; 
  signal sig000001f1 : STD_LOGIC; 
  signal sig000001f2 : STD_LOGIC; 
  signal sig000001f3 : STD_LOGIC; 
  signal sig000001f4 : STD_LOGIC; 
  signal sig000001f5 : STD_LOGIC; 
  signal sig000001f6 : STD_LOGIC; 
  signal sig000001f7 : STD_LOGIC; 
  signal sig000001f8 : STD_LOGIC; 
  signal sig000001f9 : STD_LOGIC; 
  signal sig000001fa : STD_LOGIC; 
  signal sig000001fb : STD_LOGIC; 
  signal sig000001fc : STD_LOGIC; 
  signal sig000001fd : STD_LOGIC; 
  signal sig000001fe : STD_LOGIC; 
  signal sig000001ff : STD_LOGIC; 
  signal sig00000200 : STD_LOGIC; 
  signal sig00000201 : STD_LOGIC; 
  signal sig00000202 : STD_LOGIC; 
  signal sig00000203 : STD_LOGIC; 
  signal sig00000204 : STD_LOGIC; 
  signal sig00000205 : STD_LOGIC; 
  signal sig00000206 : STD_LOGIC; 
  signal sig00000207 : STD_LOGIC; 
  signal sig00000208 : STD_LOGIC; 
  signal sig00000209 : STD_LOGIC; 
  signal sig0000020a : STD_LOGIC; 
  signal sig0000020b : STD_LOGIC; 
  signal sig0000020c : STD_LOGIC; 
  signal sig0000020d : STD_LOGIC; 
  signal sig0000020e : STD_LOGIC; 
  signal sig0000020f : STD_LOGIC; 
  signal sig00000210 : STD_LOGIC; 
  signal sig00000211 : STD_LOGIC; 
  signal sig00000212 : STD_LOGIC; 
  signal sig00000213 : STD_LOGIC; 
  signal sig00000214 : STD_LOGIC; 
  signal sig00000215 : STD_LOGIC; 
  signal sig00000216 : STD_LOGIC; 
  signal sig00000217 : STD_LOGIC; 
  signal sig00000218 : STD_LOGIC; 
  signal sig00000219 : STD_LOGIC; 
  signal sig0000021a : STD_LOGIC; 
  signal sig0000021b : STD_LOGIC; 
  signal sig0000021c : STD_LOGIC; 
  signal sig0000021d : STD_LOGIC; 
  signal sig0000021e : STD_LOGIC; 
  signal sig0000021f : STD_LOGIC; 
  signal sig00000220 : STD_LOGIC; 
  signal sig00000221 : STD_LOGIC; 
  signal sig00000222 : STD_LOGIC; 
  signal sig00000223 : STD_LOGIC; 
  signal sig00000224 : STD_LOGIC; 
  signal sig00000225 : STD_LOGIC; 
  signal sig00000226 : STD_LOGIC; 
  signal sig00000227 : STD_LOGIC; 
  signal sig00000228 : STD_LOGIC; 
  signal sig00000229 : STD_LOGIC; 
  signal sig0000022a : STD_LOGIC; 
  signal sig0000022b : STD_LOGIC; 
  signal sig0000022c : STD_LOGIC; 
  signal sig0000022d : STD_LOGIC; 
  signal sig0000022e : STD_LOGIC; 
  signal sig0000022f : STD_LOGIC; 
  signal sig00000230 : STD_LOGIC; 
  signal sig00000231 : STD_LOGIC; 
  signal sig00000232 : STD_LOGIC; 
  signal sig00000233 : STD_LOGIC; 
  signal sig00000234 : STD_LOGIC; 
  signal sig00000235 : STD_LOGIC; 
  signal sig00000236 : STD_LOGIC; 
  signal sig00000237 : STD_LOGIC; 
  signal sig00000238 : STD_LOGIC; 
  signal sig00000239 : STD_LOGIC; 
  signal sig0000023a : STD_LOGIC; 
  signal sig0000023b : STD_LOGIC; 
  signal sig0000023c : STD_LOGIC; 
  signal sig0000023d : STD_LOGIC; 
  signal sig0000023e : STD_LOGIC; 
  signal sig0000023f : STD_LOGIC; 
  signal sig00000240 : STD_LOGIC; 
  signal sig00000241 : STD_LOGIC; 
  signal sig00000242 : STD_LOGIC; 
  signal sig00000243 : STD_LOGIC; 
  signal sig00000244 : STD_LOGIC; 
  signal sig00000245 : STD_LOGIC; 
  signal sig00000246 : STD_LOGIC; 
  signal sig00000247 : STD_LOGIC; 
  signal sig00000248 : STD_LOGIC; 
  signal sig00000249 : STD_LOGIC; 
  signal sig0000024a : STD_LOGIC; 
  signal sig0000024b : STD_LOGIC; 
  signal sig0000024c : STD_LOGIC; 
  signal sig0000024d : STD_LOGIC; 
  signal sig0000024e : STD_LOGIC; 
  signal sig0000024f : STD_LOGIC; 
  signal sig00000250 : STD_LOGIC; 
  signal sig00000251 : STD_LOGIC; 
  signal sig00000252 : STD_LOGIC; 
  signal sig00000253 : STD_LOGIC; 
  signal sig00000254 : STD_LOGIC; 
  signal sig00000255 : STD_LOGIC; 
  signal sig00000256 : STD_LOGIC; 
  signal sig00000257 : STD_LOGIC; 
  signal sig00000258 : STD_LOGIC; 
  signal sig00000259 : STD_LOGIC; 
  signal sig0000025a : STD_LOGIC; 
  signal sig0000025b : STD_LOGIC; 
  signal sig0000025c : STD_LOGIC; 
  signal sig0000025d : STD_LOGIC; 
  signal sig0000025e : STD_LOGIC; 
  signal sig0000025f : STD_LOGIC; 
  signal sig00000260 : STD_LOGIC; 
  signal sig00000261 : STD_LOGIC; 
  signal sig00000262 : STD_LOGIC; 
  signal sig00000263 : STD_LOGIC; 
  signal sig00000264 : STD_LOGIC; 
  signal sig00000265 : STD_LOGIC; 
  signal sig00000266 : STD_LOGIC; 
  signal sig00000267 : STD_LOGIC; 
  signal sig00000268 : STD_LOGIC; 
  signal sig00000269 : STD_LOGIC; 
  signal sig0000026a : STD_LOGIC; 
  signal sig0000026b : STD_LOGIC; 
  signal sig0000026c : STD_LOGIC; 
  signal sig0000026d : STD_LOGIC; 
  signal sig0000026e : STD_LOGIC; 
  signal sig0000026f : STD_LOGIC; 
  signal sig00000270 : STD_LOGIC; 
  signal sig00000271 : STD_LOGIC; 
  signal sig00000272 : STD_LOGIC; 
  signal sig00000273 : STD_LOGIC; 
  signal sig00000274 : STD_LOGIC; 
  signal sig00000275 : STD_LOGIC; 
  signal sig00000276 : STD_LOGIC; 
  signal sig00000277 : STD_LOGIC; 
  signal sig00000278 : STD_LOGIC; 
  signal sig00000279 : STD_LOGIC; 
  signal sig0000027a : STD_LOGIC; 
  signal sig0000027b : STD_LOGIC; 
  signal sig0000027c : STD_LOGIC; 
  signal sig0000027d : STD_LOGIC; 
  signal sig0000027e : STD_LOGIC; 
  signal sig0000027f : STD_LOGIC; 
  signal sig00000280 : STD_LOGIC; 
  signal sig00000281 : STD_LOGIC; 
  signal sig00000282 : STD_LOGIC; 
  signal sig00000283 : STD_LOGIC; 
  signal sig00000284 : STD_LOGIC; 
  signal sig00000285 : STD_LOGIC; 
  signal sig00000286 : STD_LOGIC; 
  signal sig00000287 : STD_LOGIC; 
  signal sig00000288 : STD_LOGIC; 
  signal sig00000289 : STD_LOGIC; 
  signal sig0000028a : STD_LOGIC; 
  signal sig0000028b : STD_LOGIC; 
  signal sig0000028c : STD_LOGIC; 
  signal sig0000028d : STD_LOGIC; 
  signal sig0000028e : STD_LOGIC; 
  signal sig0000028f : STD_LOGIC; 
  signal sig00000290 : STD_LOGIC; 
  signal sig00000291 : STD_LOGIC; 
  signal sig00000292 : STD_LOGIC; 
  signal sig00000293 : STD_LOGIC; 
  signal sig00000294 : STD_LOGIC; 
  signal sig00000295 : STD_LOGIC; 
  signal sig00000296 : STD_LOGIC; 
  signal sig00000297 : STD_LOGIC; 
  signal sig00000298 : STD_LOGIC; 
  signal sig00000299 : STD_LOGIC; 
  signal sig0000029a : STD_LOGIC; 
  signal sig0000029b : STD_LOGIC; 
  signal sig0000029c : STD_LOGIC; 
  signal sig0000029d : STD_LOGIC; 
  signal sig0000029e : STD_LOGIC; 
  signal sig0000029f : STD_LOGIC; 
  signal sig000002a0 : STD_LOGIC; 
  signal sig000002a1 : STD_LOGIC; 
  signal sig000002a2 : STD_LOGIC; 
  signal sig000002a3 : STD_LOGIC; 
  signal sig000002a4 : STD_LOGIC; 
  signal sig000002a5 : STD_LOGIC; 
  signal sig000002a6 : STD_LOGIC; 
  signal sig000002a7 : STD_LOGIC; 
  signal sig000002a8 : STD_LOGIC; 
  signal sig000002a9 : STD_LOGIC; 
  signal sig000002aa : STD_LOGIC; 
  signal sig000002ab : STD_LOGIC; 
  signal sig000002ac : STD_LOGIC; 
  signal sig000002ad : STD_LOGIC; 
  signal sig000002ae : STD_LOGIC; 
  signal sig000002af : STD_LOGIC; 
  signal sig000002b0 : STD_LOGIC; 
  signal sig000002b1 : STD_LOGIC; 
  signal sig000002b2 : STD_LOGIC; 
  signal sig000002b3 : STD_LOGIC; 
  signal sig000002b4 : STD_LOGIC; 
  signal sig000002b5 : STD_LOGIC; 
  signal sig000002b6 : STD_LOGIC; 
  signal sig000002b7 : STD_LOGIC; 
  signal sig000002b8 : STD_LOGIC; 
  signal sig000002b9 : STD_LOGIC; 
  signal sig000002ba : STD_LOGIC; 
  signal sig000002bb : STD_LOGIC; 
  signal sig000002bc : STD_LOGIC; 
  signal sig000002bd : STD_LOGIC; 
  signal sig000002be : STD_LOGIC; 
  signal sig000002bf : STD_LOGIC; 
  signal sig000002c0 : STD_LOGIC; 
  signal sig000002c1 : STD_LOGIC; 
  signal sig000002c2 : STD_LOGIC; 
  signal sig000002c3 : STD_LOGIC; 
  signal sig000002c4 : STD_LOGIC; 
  signal sig000002c5 : STD_LOGIC; 
  signal sig000002c6 : STD_LOGIC; 
  signal sig000002c7 : STD_LOGIC; 
  signal sig000002c8 : STD_LOGIC; 
  signal sig000002c9 : STD_LOGIC; 
  signal sig000002ca : STD_LOGIC; 
  signal sig000002cb : STD_LOGIC; 
  signal sig000002cc : STD_LOGIC; 
  signal sig000002cd : STD_LOGIC; 
  signal sig000002ce : STD_LOGIC; 
  signal sig000002cf : STD_LOGIC; 
  signal sig000002d0 : STD_LOGIC; 
  signal sig000002d1 : STD_LOGIC; 
  signal sig000002d2 : STD_LOGIC; 
  signal sig000002d3 : STD_LOGIC; 
  signal sig000002d4 : STD_LOGIC; 
  signal sig000002d5 : STD_LOGIC; 
  signal sig000002d6 : STD_LOGIC; 
  signal sig000002d7 : STD_LOGIC; 
  signal sig000002d8 : STD_LOGIC; 
  signal sig000002d9 : STD_LOGIC; 
  signal sig000002da : STD_LOGIC; 
  signal sig000002db : STD_LOGIC; 
  signal sig000002dc : STD_LOGIC; 
  signal sig000002dd : STD_LOGIC; 
  signal sig000002de : STD_LOGIC; 
  signal sig000002df : STD_LOGIC; 
  signal sig000002e0 : STD_LOGIC; 
  signal sig000002e1 : STD_LOGIC; 
  signal sig000002e2 : STD_LOGIC; 
  signal sig000002e3 : STD_LOGIC; 
  signal sig000002e4 : STD_LOGIC; 
  signal sig000002e5 : STD_LOGIC; 
  signal sig000002e6 : STD_LOGIC; 
  signal sig000002e7 : STD_LOGIC; 
  signal sig000002e8 : STD_LOGIC; 
  signal sig000002e9 : STD_LOGIC; 
  signal sig000002ea : STD_LOGIC; 
  signal sig000002eb : STD_LOGIC; 
  signal sig000002ec : STD_LOGIC; 
  signal sig000002ed : STD_LOGIC; 
  signal sig000002ee : STD_LOGIC; 
  signal sig000002ef : STD_LOGIC; 
  signal sig000002f0 : STD_LOGIC; 
  signal sig000002f1 : STD_LOGIC; 
  signal sig000002f2 : STD_LOGIC; 
  signal sig000002f3 : STD_LOGIC; 
  signal sig000002f4 : STD_LOGIC; 
  signal sig000002f5 : STD_LOGIC; 
  signal sig000002f6 : STD_LOGIC; 
  signal sig000002f7 : STD_LOGIC; 
  signal sig000002f8 : STD_LOGIC; 
  signal sig000002f9 : STD_LOGIC; 
  signal sig000002fa : STD_LOGIC; 
  signal sig000002fb : STD_LOGIC; 
  signal sig000002fc : STD_LOGIC; 
  signal sig000002fd : STD_LOGIC; 
  signal sig000002fe : STD_LOGIC; 
  signal sig000002ff : STD_LOGIC; 
  signal sig00000300 : STD_LOGIC; 
  signal sig00000301 : STD_LOGIC; 
  signal sig00000302 : STD_LOGIC; 
  signal sig00000303 : STD_LOGIC; 
  signal sig00000304 : STD_LOGIC; 
  signal sig00000305 : STD_LOGIC; 
  signal sig00000306 : STD_LOGIC; 
  signal sig00000307 : STD_LOGIC; 
  signal sig00000308 : STD_LOGIC; 
  signal sig00000309 : STD_LOGIC; 
  signal sig0000030a : STD_LOGIC; 
  signal sig0000030b : STD_LOGIC; 
  signal sig0000030c : STD_LOGIC; 
  signal sig0000030d : STD_LOGIC; 
  signal sig0000030e : STD_LOGIC; 
  signal sig0000030f : STD_LOGIC; 
  signal sig00000310 : STD_LOGIC; 
  signal sig00000311 : STD_LOGIC; 
  signal sig00000312 : STD_LOGIC; 
  signal sig00000313 : STD_LOGIC; 
  signal sig00000314 : STD_LOGIC; 
  signal sig00000315 : STD_LOGIC; 
  signal sig00000316 : STD_LOGIC; 
  signal sig00000317 : STD_LOGIC; 
  signal sig00000318 : STD_LOGIC; 
  signal sig00000319 : STD_LOGIC; 
  signal sig0000031a : STD_LOGIC; 
  signal sig0000031b : STD_LOGIC; 
  signal sig0000031c : STD_LOGIC; 
  signal sig0000031d : STD_LOGIC; 
  signal sig0000031e : STD_LOGIC; 
  signal sig0000031f : STD_LOGIC; 
  signal sig00000320 : STD_LOGIC; 
  signal sig00000321 : STD_LOGIC; 
  signal sig00000322 : STD_LOGIC; 
  signal sig00000323 : STD_LOGIC; 
  signal sig00000324 : STD_LOGIC; 
  signal sig00000325 : STD_LOGIC; 
  signal sig00000326 : STD_LOGIC; 
  signal sig00000327 : STD_LOGIC; 
  signal sig00000328 : STD_LOGIC; 
  signal sig00000329 : STD_LOGIC; 
  signal sig0000032a : STD_LOGIC; 
  signal sig0000032b : STD_LOGIC; 
  signal sig0000032c : STD_LOGIC; 
  signal sig0000032d : STD_LOGIC; 
  signal sig0000032e : STD_LOGIC; 
  signal sig0000032f : STD_LOGIC; 
  signal sig00000330 : STD_LOGIC; 
  signal sig00000331 : STD_LOGIC; 
  signal sig00000332 : STD_LOGIC; 
  signal sig00000333 : STD_LOGIC; 
  signal sig00000334 : STD_LOGIC; 
  signal sig00000335 : STD_LOGIC; 
  signal sig00000336 : STD_LOGIC; 
  signal sig00000337 : STD_LOGIC; 
  signal sig00000338 : STD_LOGIC; 
  signal sig00000339 : STD_LOGIC; 
  signal sig0000033a : STD_LOGIC; 
  signal sig0000033b : STD_LOGIC; 
  signal sig0000033c : STD_LOGIC; 
  signal sig0000033d : STD_LOGIC; 
  signal sig0000033e : STD_LOGIC; 
  signal sig0000033f : STD_LOGIC; 
  signal sig00000340 : STD_LOGIC; 
  signal sig00000341 : STD_LOGIC; 
  signal sig00000342 : STD_LOGIC; 
  signal sig00000343 : STD_LOGIC; 
  signal sig00000344 : STD_LOGIC; 
  signal sig00000345 : STD_LOGIC; 
  signal sig00000346 : STD_LOGIC; 
  signal sig00000347 : STD_LOGIC; 
  signal sig00000348 : STD_LOGIC; 
  signal sig00000349 : STD_LOGIC; 
  signal sig0000034a : STD_LOGIC; 
  signal sig0000034b : STD_LOGIC; 
  signal sig0000034c : STD_LOGIC; 
  signal sig0000034d : STD_LOGIC; 
  signal sig0000034e : STD_LOGIC; 
  signal sig0000034f : STD_LOGIC; 
  signal sig00000350 : STD_LOGIC; 
  signal sig00000351 : STD_LOGIC; 
  signal sig00000352 : STD_LOGIC; 
  signal sig00000353 : STD_LOGIC; 
  signal sig00000354 : STD_LOGIC; 
  signal sig00000355 : STD_LOGIC; 
  signal sig00000356 : STD_LOGIC; 
  signal sig00000357 : STD_LOGIC; 
  signal sig00000358 : STD_LOGIC; 
  signal sig00000359 : STD_LOGIC; 
  signal sig0000035a : STD_LOGIC; 
  signal sig0000035b : STD_LOGIC; 
  signal sig0000035c : STD_LOGIC; 
  signal sig0000035d : STD_LOGIC; 
  signal sig0000035e : STD_LOGIC; 
  signal sig0000035f : STD_LOGIC; 
  signal sig00000360 : STD_LOGIC; 
  signal sig00000361 : STD_LOGIC; 
  signal sig00000362 : STD_LOGIC; 
  signal sig00000363 : STD_LOGIC; 
  signal sig00000364 : STD_LOGIC; 
  signal sig00000365 : STD_LOGIC; 
  signal sig00000366 : STD_LOGIC; 
  signal sig00000367 : STD_LOGIC; 
  signal sig00000368 : STD_LOGIC; 
  signal sig00000369 : STD_LOGIC; 
  signal sig0000036a : STD_LOGIC; 
  signal sig0000036b : STD_LOGIC; 
  signal sig0000036c : STD_LOGIC; 
  signal sig0000036d : STD_LOGIC; 
  signal sig0000036e : STD_LOGIC; 
  signal sig0000036f : STD_LOGIC; 
  signal sig00000370 : STD_LOGIC; 
  signal sig00000371 : STD_LOGIC; 
  signal sig00000372 : STD_LOGIC; 
  signal sig00000373 : STD_LOGIC; 
  signal sig00000374 : STD_LOGIC; 
  signal sig00000375 : STD_LOGIC; 
  signal sig00000376 : STD_LOGIC; 
  signal sig00000377 : STD_LOGIC; 
  signal sig00000378 : STD_LOGIC; 
  signal sig00000379 : STD_LOGIC; 
  signal sig0000037a : STD_LOGIC; 
  signal sig0000037b : STD_LOGIC; 
  signal sig0000037c : STD_LOGIC; 
  signal sig0000037d : STD_LOGIC; 
  signal sig0000037e : STD_LOGIC; 
  signal sig0000037f : STD_LOGIC; 
  signal sig00000380 : STD_LOGIC; 
  signal sig00000381 : STD_LOGIC; 
  signal sig00000382 : STD_LOGIC; 
  signal sig00000383 : STD_LOGIC; 
  signal sig00000384 : STD_LOGIC; 
  signal sig00000385 : STD_LOGIC; 
  signal sig00000386 : STD_LOGIC; 
  signal sig00000387 : STD_LOGIC; 
  signal sig00000388 : STD_LOGIC; 
  signal sig00000389 : STD_LOGIC; 
  signal sig0000038a : STD_LOGIC; 
  signal sig0000038b : STD_LOGIC; 
  signal sig0000038c : STD_LOGIC; 
  signal sig0000038d : STD_LOGIC; 
  signal sig0000038e : STD_LOGIC; 
  signal sig0000038f : STD_LOGIC; 
  signal sig00000390 : STD_LOGIC; 
  signal sig00000391 : STD_LOGIC; 
  signal sig00000392 : STD_LOGIC; 
  signal sig00000393 : STD_LOGIC; 
  signal sig00000394 : STD_LOGIC; 
  signal sig00000395 : STD_LOGIC; 
  signal sig00000396 : STD_LOGIC; 
  signal sig00000397 : STD_LOGIC; 
  signal sig00000398 : STD_LOGIC; 
  signal sig00000399 : STD_LOGIC; 
  signal sig0000039a : STD_LOGIC; 
  signal sig0000039b : STD_LOGIC; 
  signal sig0000039c : STD_LOGIC; 
  signal sig0000039d : STD_LOGIC; 
  signal sig0000039e : STD_LOGIC; 
  signal sig0000039f : STD_LOGIC; 
  signal sig000003a0 : STD_LOGIC; 
  signal sig000003a1 : STD_LOGIC; 
  signal sig000003a2 : STD_LOGIC; 
  signal sig000003a3 : STD_LOGIC; 
  signal sig000003a4 : STD_LOGIC; 
  signal sig000003a5 : STD_LOGIC; 
  signal sig000003a6 : STD_LOGIC; 
  signal sig000003a7 : STD_LOGIC; 
  signal sig000003a8 : STD_LOGIC; 
  signal sig000003a9 : STD_LOGIC; 
  signal sig000003aa : STD_LOGIC; 
  signal sig000003ab : STD_LOGIC; 
  signal sig000003ac : STD_LOGIC; 
  signal sig000003ad : STD_LOGIC; 
  signal sig000003ae : STD_LOGIC; 
  signal sig000003af : STD_LOGIC; 
  signal sig000003b0 : STD_LOGIC; 
  signal sig000003b1 : STD_LOGIC; 
  signal sig000003b2 : STD_LOGIC; 
  signal sig000003b3 : STD_LOGIC; 
  signal sig000003b4 : STD_LOGIC; 
  signal sig000003b5 : STD_LOGIC; 
  signal sig000003b6 : STD_LOGIC; 
  signal sig000003b7 : STD_LOGIC; 
  signal sig000003b8 : STD_LOGIC; 
  signal sig000003b9 : STD_LOGIC; 
  signal sig000003ba : STD_LOGIC; 
  signal sig000003bb : STD_LOGIC; 
  signal sig000003bc : STD_LOGIC; 
  signal sig000003bd : STD_LOGIC; 
  signal sig000003be : STD_LOGIC; 
  signal sig000003bf : STD_LOGIC; 
  signal sig000003c0 : STD_LOGIC; 
  signal sig000003c1 : STD_LOGIC; 
  signal sig000003c2 : STD_LOGIC; 
  signal sig000003c3 : STD_LOGIC; 
  signal sig000003c4 : STD_LOGIC; 
  signal sig000003c5 : STD_LOGIC; 
  signal sig000003c6 : STD_LOGIC; 
  signal sig000003c7 : STD_LOGIC; 
  signal sig000003c8 : STD_LOGIC; 
  signal sig000003c9 : STD_LOGIC; 
  signal sig000003ca : STD_LOGIC; 
  signal sig000003cb : STD_LOGIC; 
  signal sig000003cc : STD_LOGIC; 
  signal sig000003cd : STD_LOGIC; 
  signal sig000003ce : STD_LOGIC; 
  signal sig000003cf : STD_LOGIC; 
  signal sig000003d0 : STD_LOGIC; 
  signal sig000003d1 : STD_LOGIC; 
  signal sig000003d2 : STD_LOGIC; 
  signal sig000003d3 : STD_LOGIC; 
  signal sig000003d4 : STD_LOGIC; 
  signal sig000003d5 : STD_LOGIC; 
  signal sig000003d6 : STD_LOGIC; 
  signal sig000003d7 : STD_LOGIC; 
  signal sig000003d8 : STD_LOGIC; 
  signal sig000003d9 : STD_LOGIC; 
  signal sig000003da : STD_LOGIC; 
  signal sig000003db : STD_LOGIC; 
  signal sig000003dc : STD_LOGIC; 
  signal sig000003dd : STD_LOGIC; 
  signal sig000003de : STD_LOGIC; 
  signal sig000003df : STD_LOGIC; 
  signal sig000003e0 : STD_LOGIC; 
  signal sig000003e1 : STD_LOGIC; 
  signal sig000003e2 : STD_LOGIC; 
  signal sig000003e3 : STD_LOGIC; 
  signal sig000003e4 : STD_LOGIC; 
  signal sig000003e5 : STD_LOGIC; 
  signal sig000003e6 : STD_LOGIC; 
  signal sig000003e7 : STD_LOGIC; 
  signal sig000003e8 : STD_LOGIC; 
  signal sig000003e9 : STD_LOGIC; 
  signal sig000003ea : STD_LOGIC; 
  signal sig000003eb : STD_LOGIC; 
  signal sig000003ec : STD_LOGIC; 
  signal sig000003ed : STD_LOGIC; 
  signal sig000003ee : STD_LOGIC; 
  signal sig000003ef : STD_LOGIC; 
  signal sig000003f0 : STD_LOGIC; 
  signal sig000003f1 : STD_LOGIC; 
  signal sig000003f2 : STD_LOGIC; 
  signal sig000003f3 : STD_LOGIC; 
  signal sig000003f4 : STD_LOGIC; 
  signal sig000003f5 : STD_LOGIC; 
  signal sig000003f6 : STD_LOGIC; 
  signal sig000003f7 : STD_LOGIC; 
  signal sig000003f8 : STD_LOGIC; 
  signal sig000003f9 : STD_LOGIC; 
  signal sig000003fa : STD_LOGIC; 
  signal sig000003fb : STD_LOGIC; 
  signal sig000003fc : STD_LOGIC; 
  signal sig000003fd : STD_LOGIC; 
  signal sig000003fe : STD_LOGIC; 
  signal sig000003ff : STD_LOGIC; 
  signal sig00000400 : STD_LOGIC; 
  signal sig00000401 : STD_LOGIC; 
  signal sig00000402 : STD_LOGIC; 
  signal sig00000403 : STD_LOGIC; 
  signal sig00000404 : STD_LOGIC; 
  signal sig00000405 : STD_LOGIC; 
  signal sig00000406 : STD_LOGIC; 
  signal sig00000407 : STD_LOGIC; 
  signal sig00000408 : STD_LOGIC; 
  signal sig00000409 : STD_LOGIC; 
  signal sig0000040a : STD_LOGIC; 
  signal sig0000040b : STD_LOGIC; 
  signal sig0000040c : STD_LOGIC; 
  signal sig0000040d : STD_LOGIC; 
  signal sig0000040e : STD_LOGIC; 
  signal sig0000040f : STD_LOGIC; 
  signal sig00000410 : STD_LOGIC; 
  signal sig00000411 : STD_LOGIC; 
  signal sig00000412 : STD_LOGIC; 
  signal sig00000413 : STD_LOGIC; 
  signal sig00000414 : STD_LOGIC; 
  signal sig00000415 : STD_LOGIC; 
  signal sig00000416 : STD_LOGIC; 
  signal sig00000417 : STD_LOGIC; 
  signal sig00000418 : STD_LOGIC; 
  signal sig00000419 : STD_LOGIC; 
  signal sig0000041a : STD_LOGIC; 
  signal sig0000041b : STD_LOGIC; 
  signal sig0000041c : STD_LOGIC; 
  signal sig0000041d : STD_LOGIC; 
  signal sig0000041e : STD_LOGIC; 
  signal sig0000041f : STD_LOGIC; 
  signal sig00000420 : STD_LOGIC; 
  signal sig00000421 : STD_LOGIC; 
  signal sig00000422 : STD_LOGIC; 
  signal sig00000423 : STD_LOGIC; 
  signal sig00000424 : STD_LOGIC; 
  signal sig00000425 : STD_LOGIC; 
  signal sig00000426 : STD_LOGIC; 
  signal sig00000427 : STD_LOGIC; 
  signal sig00000428 : STD_LOGIC; 
  signal sig00000429 : STD_LOGIC; 
  signal sig0000042a : STD_LOGIC; 
  signal sig0000042b : STD_LOGIC; 
  signal sig0000042c : STD_LOGIC; 
  signal sig0000042d : STD_LOGIC; 
  signal sig0000042e : STD_LOGIC; 
  signal sig0000042f : STD_LOGIC; 
  signal sig00000430 : STD_LOGIC; 
  signal sig00000431 : STD_LOGIC; 
  signal sig00000432 : STD_LOGIC; 
  signal sig00000433 : STD_LOGIC; 
  signal sig00000434 : STD_LOGIC; 
  signal sig00000435 : STD_LOGIC; 
  signal sig00000436 : STD_LOGIC; 
  signal sig00000437 : STD_LOGIC; 
  signal sig00000438 : STD_LOGIC; 
  signal sig00000439 : STD_LOGIC; 
  signal sig0000043a : STD_LOGIC; 
  signal sig0000043b : STD_LOGIC; 
  signal sig0000043c : STD_LOGIC; 
  signal sig0000043d : STD_LOGIC; 
  signal sig0000043e : STD_LOGIC; 
  signal sig0000043f : STD_LOGIC; 
  signal sig00000440 : STD_LOGIC; 
  signal sig00000441 : STD_LOGIC; 
  signal sig00000442 : STD_LOGIC; 
  signal sig00000443 : STD_LOGIC; 
  signal sig00000444 : STD_LOGIC; 
  signal sig00000445 : STD_LOGIC; 
  signal sig00000446 : STD_LOGIC; 
  signal sig00000447 : STD_LOGIC; 
  signal sig00000448 : STD_LOGIC; 
  signal sig00000449 : STD_LOGIC; 
  signal sig0000044a : STD_LOGIC; 
  signal sig0000044b : STD_LOGIC; 
  signal sig0000044c : STD_LOGIC; 
  signal sig0000044d : STD_LOGIC; 
  signal sig0000044e : STD_LOGIC; 
  signal sig0000044f : STD_LOGIC; 
  signal sig00000450 : STD_LOGIC; 
  signal sig00000451 : STD_LOGIC; 
  signal sig00000452 : STD_LOGIC; 
  signal sig00000453 : STD_LOGIC; 
  signal sig00000454 : STD_LOGIC; 
  signal sig00000455 : STD_LOGIC; 
  signal sig00000456 : STD_LOGIC; 
  signal sig00000457 : STD_LOGIC; 
  signal sig00000458 : STD_LOGIC; 
  signal sig00000459 : STD_LOGIC; 
  signal sig0000045a : STD_LOGIC; 
  signal sig0000045b : STD_LOGIC; 
  signal sig0000045c : STD_LOGIC; 
  signal sig0000045d : STD_LOGIC; 
  signal sig0000045e : STD_LOGIC; 
  signal sig0000045f : STD_LOGIC; 
  signal sig00000460 : STD_LOGIC; 
  signal sig00000461 : STD_LOGIC; 
  signal sig00000462 : STD_LOGIC; 
  signal sig00000463 : STD_LOGIC; 
  signal sig00000464 : STD_LOGIC; 
  signal sig00000465 : STD_LOGIC; 
  signal sig00000466 : STD_LOGIC; 
  signal sig00000467 : STD_LOGIC; 
  signal sig00000468 : STD_LOGIC; 
  signal sig00000469 : STD_LOGIC; 
  signal sig0000046a : STD_LOGIC; 
  signal sig0000046b : STD_LOGIC; 
  signal sig0000046c : STD_LOGIC; 
  signal sig0000046d : STD_LOGIC; 
  signal sig0000046e : STD_LOGIC; 
  signal sig0000046f : STD_LOGIC; 
  signal sig00000470 : STD_LOGIC; 
  signal sig00000471 : STD_LOGIC; 
  signal sig00000472 : STD_LOGIC; 
  signal sig00000473 : STD_LOGIC; 
  signal sig00000474 : STD_LOGIC; 
  signal sig00000475 : STD_LOGIC; 
  signal sig00000476 : STD_LOGIC; 
  signal sig00000477 : STD_LOGIC; 
  signal sig00000478 : STD_LOGIC; 
  signal sig00000479 : STD_LOGIC; 
  signal sig0000047a : STD_LOGIC; 
  signal sig0000047b : STD_LOGIC; 
  signal sig0000047c : STD_LOGIC; 
  signal sig0000047d : STD_LOGIC; 
  signal sig0000047e : STD_LOGIC; 
  signal sig0000047f : STD_LOGIC; 
  signal sig00000480 : STD_LOGIC; 
  signal sig00000481 : STD_LOGIC; 
  signal sig00000482 : STD_LOGIC; 
  signal sig00000483 : STD_LOGIC; 
  signal sig00000484 : STD_LOGIC; 
  signal sig00000485 : STD_LOGIC; 
  signal sig00000486 : STD_LOGIC; 
  signal sig00000487 : STD_LOGIC; 
  signal sig00000488 : STD_LOGIC; 
  signal sig00000489 : STD_LOGIC; 
  signal sig0000048a : STD_LOGIC; 
  signal sig0000048b : STD_LOGIC; 
  signal sig0000048c : STD_LOGIC; 
  signal sig0000048d : STD_LOGIC; 
  signal sig0000048e : STD_LOGIC; 
  signal sig0000048f : STD_LOGIC; 
  signal sig00000490 : STD_LOGIC; 
  signal sig00000491 : STD_LOGIC; 
  signal sig00000492 : STD_LOGIC; 
  signal sig00000493 : STD_LOGIC; 
  signal sig00000494 : STD_LOGIC; 
  signal sig00000495 : STD_LOGIC; 
  signal sig00000496 : STD_LOGIC; 
  signal sig00000497 : STD_LOGIC; 
  signal sig00000498 : STD_LOGIC; 
  signal sig00000499 : STD_LOGIC; 
  signal sig0000049a : STD_LOGIC; 
  signal sig0000049b : STD_LOGIC; 
  signal sig0000049c : STD_LOGIC; 
  signal sig0000049d : STD_LOGIC; 
  signal sig0000049e : STD_LOGIC; 
  signal sig0000049f : STD_LOGIC; 
  signal sig000004a0 : STD_LOGIC; 
  signal sig000004a1 : STD_LOGIC; 
  signal sig000004a2 : STD_LOGIC; 
  signal sig000004a3 : STD_LOGIC; 
  signal sig000004a4 : STD_LOGIC; 
  signal sig000004a5 : STD_LOGIC; 
  signal sig000004a6 : STD_LOGIC; 
  signal sig000004a7 : STD_LOGIC; 
  signal sig000004a8 : STD_LOGIC; 
  signal sig000004a9 : STD_LOGIC; 
  signal sig000004aa : STD_LOGIC; 
  signal sig000004ab : STD_LOGIC; 
  signal sig000004ac : STD_LOGIC; 
  signal sig000004ad : STD_LOGIC; 
  signal sig000004ae : STD_LOGIC; 
  signal sig000004af : STD_LOGIC; 
  signal sig000004b0 : STD_LOGIC; 
  signal sig000004b1 : STD_LOGIC; 
  signal sig000004b2 : STD_LOGIC; 
  signal sig000004b3 : STD_LOGIC; 
  signal sig000004b4 : STD_LOGIC; 
  signal sig000004b5 : STD_LOGIC; 
  signal sig000004b6 : STD_LOGIC; 
  signal sig000004b7 : STD_LOGIC; 
  signal sig000004b8 : STD_LOGIC; 
  signal sig000004b9 : STD_LOGIC; 
  signal sig000004ba : STD_LOGIC; 
  signal sig000004bb : STD_LOGIC; 
  signal sig000004bc : STD_LOGIC; 
  signal sig000004bd : STD_LOGIC; 
  signal sig000004be : STD_LOGIC; 
  signal sig000004bf : STD_LOGIC; 
  signal sig000004c0 : STD_LOGIC; 
  signal sig000004c1 : STD_LOGIC; 
  signal sig000004c2 : STD_LOGIC; 
  signal sig000004c3 : STD_LOGIC; 
  signal sig000004c4 : STD_LOGIC; 
  signal sig000004c5 : STD_LOGIC; 
  signal sig000004c6 : STD_LOGIC; 
  signal sig000004c7 : STD_LOGIC; 
  signal sig000004c8 : STD_LOGIC; 
  signal sig000004c9 : STD_LOGIC; 
  signal sig000004ca : STD_LOGIC; 
  signal sig000004cb : STD_LOGIC; 
  signal sig000004cc : STD_LOGIC; 
  signal sig000004cd : STD_LOGIC; 
  signal sig000004ce : STD_LOGIC; 
  signal sig000004cf : STD_LOGIC; 
  signal sig000004d0 : STD_LOGIC; 
  signal sig000004d1 : STD_LOGIC; 
  signal sig000004d2 : STD_LOGIC; 
  signal sig000004d3 : STD_LOGIC; 
  signal sig000004d4 : STD_LOGIC; 
  signal sig000004d5 : STD_LOGIC; 
  signal sig000004d6 : STD_LOGIC; 
  signal sig000004d7 : STD_LOGIC; 
  signal sig000004d8 : STD_LOGIC; 
  signal sig000004d9 : STD_LOGIC; 
  signal sig000004da : STD_LOGIC; 
  signal sig000004db : STD_LOGIC; 
  signal sig000004dc : STD_LOGIC; 
  signal sig000004dd : STD_LOGIC; 
  signal sig000004de : STD_LOGIC; 
  signal sig000004df : STD_LOGIC; 
  signal sig000004e0 : STD_LOGIC; 
  signal sig000004e1 : STD_LOGIC; 
  signal sig000004e2 : STD_LOGIC; 
  signal sig000004e3 : STD_LOGIC; 
  signal sig000004e4 : STD_LOGIC; 
  signal sig000004e5 : STD_LOGIC; 
  signal sig000004e6 : STD_LOGIC; 
  signal sig000004e7 : STD_LOGIC; 
  signal sig000004e8 : STD_LOGIC; 
  signal sig000004e9 : STD_LOGIC; 
  signal sig000004ea : STD_LOGIC; 
  signal sig000004eb : STD_LOGIC; 
  signal sig000004ec : STD_LOGIC; 
  signal sig000004ed : STD_LOGIC; 
  signal sig000004ee : STD_LOGIC; 
  signal sig000004ef : STD_LOGIC; 
  signal sig000004f0 : STD_LOGIC; 
  signal sig000004f1 : STD_LOGIC; 
  signal sig000004f2 : STD_LOGIC; 
  signal sig000004f3 : STD_LOGIC; 
  signal sig000004f4 : STD_LOGIC; 
  signal sig000004f5 : STD_LOGIC; 
  signal sig000004f6 : STD_LOGIC; 
  signal sig000004f7 : STD_LOGIC; 
  signal sig000004f8 : STD_LOGIC; 
  signal sig000004f9 : STD_LOGIC; 
  signal sig000004fa : STD_LOGIC; 
  signal sig000004fb : STD_LOGIC; 
  signal sig000004fc : STD_LOGIC; 
  signal sig000004fd : STD_LOGIC; 
  signal sig000004fe : STD_LOGIC; 
  signal sig000004ff : STD_LOGIC; 
  signal sig00000500 : STD_LOGIC; 
  signal sig00000501 : STD_LOGIC; 
  signal sig00000502 : STD_LOGIC; 
  signal sig00000503 : STD_LOGIC; 
  signal sig00000504 : STD_LOGIC; 
  signal sig00000505 : STD_LOGIC; 
  signal sig00000506 : STD_LOGIC; 
  signal sig00000507 : STD_LOGIC; 
  signal sig00000508 : STD_LOGIC; 
  signal sig00000509 : STD_LOGIC; 
  signal sig0000050a : STD_LOGIC; 
  signal sig0000050b : STD_LOGIC; 
  signal sig0000050c : STD_LOGIC; 
  signal sig0000050d : STD_LOGIC; 
  signal sig0000050e : STD_LOGIC; 
  signal sig0000050f : STD_LOGIC; 
  signal sig00000510 : STD_LOGIC; 
  signal sig00000511 : STD_LOGIC; 
  signal sig00000512 : STD_LOGIC; 
  signal sig00000513 : STD_LOGIC; 
  signal sig00000514 : STD_LOGIC; 
  signal sig00000515 : STD_LOGIC; 
  signal sig0000052a : STD_LOGIC; 
  signal sig0000052b : STD_LOGIC; 
  signal sig0000052c : STD_LOGIC; 
  signal sig0000052d : STD_LOGIC; 
  signal sig0000052e : STD_LOGIC; 
  signal sig0000052f : STD_LOGIC; 
  signal sig00000530 : STD_LOGIC; 
  signal sig0000053d : STD_LOGIC; 
  signal sig0000053e : STD_LOGIC; 
  signal sig0000053f : STD_LOGIC; 
  signal sig00000540 : STD_LOGIC; 
  signal sig00000541 : STD_LOGIC; 
  signal sig00000542 : STD_LOGIC; 
  signal sig00000543 : STD_LOGIC; 
  signal sig00000544 : STD_LOGIC; 
  signal sig00000545 : STD_LOGIC; 
  signal sig00000546 : STD_LOGIC; 
  signal sig00000547 : STD_LOGIC; 
  signal sig00000548 : STD_LOGIC; 
  signal sig00000549 : STD_LOGIC; 
  signal sig0000054d : STD_LOGIC; 
  signal sig0000054e : STD_LOGIC; 
  signal sig0000054f : STD_LOGIC; 
  signal sig00000550 : STD_LOGIC; 
  signal sig00000551 : STD_LOGIC; 
  signal sig00000552 : STD_LOGIC; 
  signal sig00000553 : STD_LOGIC; 
  signal sig00000554 : STD_LOGIC; 
  signal sig00000555 : STD_LOGIC; 
  signal sig00000556 : STD_LOGIC; 
  signal sig00000557 : STD_LOGIC; 
  signal sig00000558 : STD_LOGIC; 
  signal sig00000559 : STD_LOGIC; 
  signal sig0000055a : STD_LOGIC; 
  signal sig0000055b : STD_LOGIC; 
  signal sig0000055c : STD_LOGIC; 
  signal sig0000055d : STD_LOGIC; 
  signal sig0000055e : STD_LOGIC; 
  signal sig0000055f : STD_LOGIC; 
  signal sig00000560 : STD_LOGIC; 
  signal sig00000561 : STD_LOGIC; 
  signal sig00000562 : STD_LOGIC; 
  signal sig00000563 : STD_LOGIC; 
  signal sig00000564 : STD_LOGIC; 
  signal sig00000565 : STD_LOGIC; 
  signal sig00000566 : STD_LOGIC; 
  signal sig00000567 : STD_LOGIC; 
  signal sig00000568 : STD_LOGIC; 
  signal sig00000569 : STD_LOGIC; 
  signal sig0000056a : STD_LOGIC; 
  signal sig0000056b : STD_LOGIC; 
  signal sig0000056c : STD_LOGIC; 
  signal sig0000056d : STD_LOGIC; 
  signal sig0000056e : STD_LOGIC; 
  signal sig0000056f : STD_LOGIC; 
  signal sig00000570 : STD_LOGIC; 
  signal sig00000571 : STD_LOGIC; 
  signal sig00000572 : STD_LOGIC; 
  signal sig00000573 : STD_LOGIC; 
  signal sig00000574 : STD_LOGIC; 
  signal sig00000575 : STD_LOGIC; 
  signal sig00000576 : STD_LOGIC; 
  signal sig00000577 : STD_LOGIC; 
  signal sig00000578 : STD_LOGIC; 
  signal sig00000579 : STD_LOGIC; 
  signal sig0000057a : STD_LOGIC; 
  signal sig0000057b : STD_LOGIC; 
  signal sig0000057c : STD_LOGIC; 
  signal sig0000057d : STD_LOGIC; 
  signal sig0000057e : STD_LOGIC; 
  signal sig0000057f : STD_LOGIC; 
  signal sig00000580 : STD_LOGIC; 
  signal sig00000581 : STD_LOGIC; 
  signal sig00000582 : STD_LOGIC; 
  signal sig00000583 : STD_LOGIC; 
  signal sig00000584 : STD_LOGIC; 
  signal sig00000585 : STD_LOGIC; 
  signal sig00000586 : STD_LOGIC; 
  signal sig00000592 : STD_LOGIC; 
  signal sig00000593 : STD_LOGIC; 
  signal sig00000594 : STD_LOGIC; 
  signal sig00000595 : STD_LOGIC; 
  signal sig00000596 : STD_LOGIC; 
  signal sig00000597 : STD_LOGIC; 
  signal sig00000598 : STD_LOGIC; 
  signal sig00000599 : STD_LOGIC; 
  signal sig0000059a : STD_LOGIC; 
  signal sig0000059b : STD_LOGIC; 
  signal sig0000059c : STD_LOGIC; 
  signal sig0000059d : STD_LOGIC; 
  signal sig0000059e : STD_LOGIC; 
  signal sig0000059f : STD_LOGIC; 
  signal sig000005a4 : STD_LOGIC; 
  signal sig000005a5 : STD_LOGIC; 
  signal sig000005a6 : STD_LOGIC; 
  signal sig000005a7 : STD_LOGIC; 
  signal sig000005a8 : STD_LOGIC; 
  signal sig000005a9 : STD_LOGIC; 
  signal sig000005aa : STD_LOGIC; 
  signal sig000005ab : STD_LOGIC; 
  signal sig000005ac : STD_LOGIC; 
  signal sig000005ad : STD_LOGIC; 
  signal sig000005ae : STD_LOGIC; 
  signal sig000005af : STD_LOGIC; 
  signal sig000005b0 : STD_LOGIC; 
  signal sig000005b1 : STD_LOGIC; 
  signal sig000005b2 : STD_LOGIC; 
  signal sig000005b3 : STD_LOGIC; 
  signal sig000005b4 : STD_LOGIC; 
  signal sig000005b5 : STD_LOGIC; 
  signal sig000005b6 : STD_LOGIC; 
  signal sig000005b7 : STD_LOGIC; 
  signal sig000005b8 : STD_LOGIC; 
  signal sig000005b9 : STD_LOGIC; 
  signal sig000005ba : STD_LOGIC; 
  signal sig000005bb : STD_LOGIC; 
  signal sig000005bc : STD_LOGIC; 
  signal sig000005bd : STD_LOGIC; 
  signal sig000005be : STD_LOGIC; 
  signal sig000005bf : STD_LOGIC; 
  signal sig000005c0 : STD_LOGIC; 
  signal sig000005c1 : STD_LOGIC; 
  signal sig000005d6 : STD_LOGIC; 
  signal sig000005d7 : STD_LOGIC; 
  signal sig000005d8 : STD_LOGIC; 
  signal sig000005d9 : STD_LOGIC; 
  signal sig000005da : STD_LOGIC; 
  signal sig000005db : STD_LOGIC; 
  signal sig000005dc : STD_LOGIC; 
  signal sig000005e9 : STD_LOGIC; 
  signal sig000005ea : STD_LOGIC; 
  signal sig000005eb : STD_LOGIC; 
  signal sig000005ec : STD_LOGIC; 
  signal sig000005ed : STD_LOGIC; 
  signal sig000005ee : STD_LOGIC; 
  signal sig000005ef : STD_LOGIC; 
  signal sig000005f0 : STD_LOGIC; 
  signal sig000005f1 : STD_LOGIC; 
  signal sig000005f2 : STD_LOGIC; 
  signal sig000005f3 : STD_LOGIC; 
  signal sig000005f4 : STD_LOGIC; 
  signal sig000005f5 : STD_LOGIC; 
  signal sig000005f9 : STD_LOGIC; 
  signal sig000005fa : STD_LOGIC; 
  signal sig000005fb : STD_LOGIC; 
  signal sig000005fc : STD_LOGIC; 
  signal sig000005fd : STD_LOGIC; 
  signal sig000005fe : STD_LOGIC; 
  signal sig000005ff : STD_LOGIC; 
  signal sig00000600 : STD_LOGIC; 
  signal sig00000601 : STD_LOGIC; 
  signal sig00000602 : STD_LOGIC; 
  signal sig00000603 : STD_LOGIC; 
  signal sig00000604 : STD_LOGIC; 
  signal sig00000605 : STD_LOGIC; 
  signal sig00000607 : STD_LOGIC; 
  signal sig00000608 : STD_LOGIC; 
  signal sig00000609 : STD_LOGIC; 
  signal sig0000060a : STD_LOGIC; 
  signal sig0000060b : STD_LOGIC; 
  signal sig0000060c : STD_LOGIC; 
  signal sig0000060d : STD_LOGIC; 
  signal sig0000060e : STD_LOGIC; 
  signal sig0000060f : STD_LOGIC; 
  signal sig00000610 : STD_LOGIC; 
  signal sig00000611 : STD_LOGIC; 
  signal sig00000612 : STD_LOGIC; 
  signal sig00000613 : STD_LOGIC; 
  signal sig00000614 : STD_LOGIC; 
  signal sig00000615 : STD_LOGIC; 
  signal sig00000616 : STD_LOGIC; 
  signal sig00000617 : STD_LOGIC; 
  signal sig00000618 : STD_LOGIC; 
  signal sig00000619 : STD_LOGIC; 
  signal sig0000061a : STD_LOGIC; 
  signal sig0000061b : STD_LOGIC; 
  signal sig0000061c : STD_LOGIC; 
  signal sig0000061d : STD_LOGIC; 
  signal sig0000061e : STD_LOGIC; 
  signal sig0000061f : STD_LOGIC; 
  signal sig00000620 : STD_LOGIC; 
  signal sig00000621 : STD_LOGIC; 
  signal sig00000622 : STD_LOGIC; 
  signal sig00000623 : STD_LOGIC; 
  signal sig00000624 : STD_LOGIC; 
  signal sig00000625 : STD_LOGIC; 
  signal sig00000626 : STD_LOGIC; 
  signal sig00000627 : STD_LOGIC; 
  signal sig00000628 : STD_LOGIC; 
  signal sig00000629 : STD_LOGIC; 
  signal sig0000062a : STD_LOGIC; 
  signal sig0000062b : STD_LOGIC; 
  signal sig0000062c : STD_LOGIC; 
  signal sig0000062d : STD_LOGIC; 
  signal sig0000062e : STD_LOGIC; 
  signal sig0000062f : STD_LOGIC; 
  signal sig00000630 : STD_LOGIC; 
  signal sig00000631 : STD_LOGIC; 
  signal sig00000632 : STD_LOGIC; 
  signal sig00000633 : STD_LOGIC; 
  signal sig00000634 : STD_LOGIC; 
  signal sig00000635 : STD_LOGIC; 
  signal sig00000636 : STD_LOGIC; 
  signal sig00000637 : STD_LOGIC; 
  signal sig00000638 : STD_LOGIC; 
  signal sig00000639 : STD_LOGIC; 
  signal sig000006a9 : STD_LOGIC; 
  signal sig000006aa : STD_LOGIC; 
  signal sig000006ab : STD_LOGIC; 
  signal sig000006ac : STD_LOGIC; 
  signal sig000006ad : STD_LOGIC; 
  signal sig000006ae : STD_LOGIC; 
  signal sig000006af : STD_LOGIC; 
  signal sig000006b0 : STD_LOGIC; 
  signal sig000006b1 : STD_LOGIC; 
  signal sig000006b2 : STD_LOGIC; 
  signal sig000006b3 : STD_LOGIC; 
  signal sig000006b4 : STD_LOGIC; 
  signal sig000006b5 : STD_LOGIC; 
  signal sig000006b6 : STD_LOGIC; 
  signal sig000006b7 : STD_LOGIC; 
  signal sig000006b8 : STD_LOGIC; 
  signal sig000006b9 : STD_LOGIC; 
  signal sig000006ba : STD_LOGIC; 
  signal sig000006bb : STD_LOGIC; 
  signal sig000006bc : STD_LOGIC; 
  signal sig000006bd : STD_LOGIC; 
  signal sig000006be : STD_LOGIC; 
  signal sig000006bf : STD_LOGIC; 
  signal sig000006c0 : STD_LOGIC; 
  signal sig000006c1 : STD_LOGIC; 
  signal sig000006c2 : STD_LOGIC; 
  signal sig000006c3 : STD_LOGIC; 
  signal sig000006c4 : STD_LOGIC; 
  signal sig000006c5 : STD_LOGIC; 
  signal sig000006c6 : STD_LOGIC; 
  signal sig000006c7 : STD_LOGIC; 
  signal sig000006c8 : STD_LOGIC; 
  signal sig000006c9 : STD_LOGIC; 
  signal sig000006ca : STD_LOGIC; 
  signal sig000006cb : STD_LOGIC; 
  signal sig000006cc : STD_LOGIC; 
  signal sig000006cd : STD_LOGIC; 
  signal sig000006ce : STD_LOGIC; 
  signal sig000006cf : STD_LOGIC; 
  signal sig000006d0 : STD_LOGIC; 
  signal sig000006d1 : STD_LOGIC; 
  signal sig000006d2 : STD_LOGIC; 
  signal sig000006d3 : STD_LOGIC; 
  signal sig000006d4 : STD_LOGIC; 
  signal sig000006d5 : STD_LOGIC; 
  signal sig000006d6 : STD_LOGIC; 
  signal sig000006d7 : STD_LOGIC; 
  signal sig000006d8 : STD_LOGIC; 
  signal sig000006d9 : STD_LOGIC; 
  signal sig000006da : STD_LOGIC; 
  signal sig000006db : STD_LOGIC; 
  signal sig000006dc : STD_LOGIC; 
  signal sig000006dd : STD_LOGIC; 
  signal sig000006de : STD_LOGIC; 
  signal sig000006df : STD_LOGIC; 
  signal sig000006e0 : STD_LOGIC; 
  signal sig000006e1 : STD_LOGIC; 
  signal sig000006e2 : STD_LOGIC; 
  signal sig000006e3 : STD_LOGIC; 
  signal sig000006e4 : STD_LOGIC; 
  signal sig000006e5 : STD_LOGIC; 
  signal sig000006e6 : STD_LOGIC; 
  signal sig000006e7 : STD_LOGIC; 
  signal sig000006e8 : STD_LOGIC; 
  signal sig000006e9 : STD_LOGIC; 
  signal sig000006ea : STD_LOGIC; 
  signal sig000006eb : STD_LOGIC; 
  signal sig000006ec : STD_LOGIC; 
  signal sig000006ed : STD_LOGIC; 
  signal sig000006ee : STD_LOGIC; 
  signal sig000006ef : STD_LOGIC; 
  signal sig000006f0 : STD_LOGIC; 
  signal sig000006f1 : STD_LOGIC; 
  signal sig000006f2 : STD_LOGIC; 
  signal sig000006f3 : STD_LOGIC; 
  signal sig000006f4 : STD_LOGIC; 
  signal sig000006f5 : STD_LOGIC; 
  signal sig000006f6 : STD_LOGIC; 
  signal sig000006f7 : STD_LOGIC; 
  signal sig000006f8 : STD_LOGIC; 
  signal sig000006f9 : STD_LOGIC; 
  signal sig000006fa : STD_LOGIC; 
  signal sig000006fb : STD_LOGIC; 
  signal sig000006fc : STD_LOGIC; 
  signal sig000006fd : STD_LOGIC; 
  signal sig000006fe : STD_LOGIC; 
  signal sig000006ff : STD_LOGIC; 
  signal sig00000700 : STD_LOGIC; 
  signal sig00000701 : STD_LOGIC; 
  signal sig00000702 : STD_LOGIC; 
  signal sig00000703 : STD_LOGIC; 
  signal sig00000704 : STD_LOGIC; 
  signal sig00000705 : STD_LOGIC; 
  signal sig00000706 : STD_LOGIC; 
  signal sig00000707 : STD_LOGIC; 
  signal sig00000708 : STD_LOGIC; 
  signal sig00000709 : STD_LOGIC; 
  signal sig0000070a : STD_LOGIC; 
  signal sig0000070b : STD_LOGIC; 
  signal sig0000070c : STD_LOGIC; 
  signal sig0000070d : STD_LOGIC; 
  signal sig0000070e : STD_LOGIC; 
  signal sig0000070f : STD_LOGIC; 
  signal sig00000710 : STD_LOGIC; 
  signal sig00000711 : STD_LOGIC; 
  signal sig00000712 : STD_LOGIC; 
  signal sig00000713 : STD_LOGIC; 
  signal sig00000714 : STD_LOGIC; 
  signal sig00000715 : STD_LOGIC; 
  signal sig00000716 : STD_LOGIC; 
  signal sig00000717 : STD_LOGIC; 
  signal sig00000718 : STD_LOGIC; 
  signal sig00000719 : STD_LOGIC; 
  signal sig0000071a : STD_LOGIC; 
  signal sig0000071b : STD_LOGIC; 
  signal sig0000071c : STD_LOGIC; 
  signal sig0000071d : STD_LOGIC; 
  signal sig0000071e : STD_LOGIC; 
  signal sig0000071f : STD_LOGIC; 
  signal sig00000720 : STD_LOGIC; 
  signal sig00000721 : STD_LOGIC; 
  signal sig00000722 : STD_LOGIC; 
  signal sig00000723 : STD_LOGIC; 
  signal sig00000724 : STD_LOGIC; 
  signal sig00000725 : STD_LOGIC; 
  signal sig00000726 : STD_LOGIC; 
  signal sig00000727 : STD_LOGIC; 
  signal sig00000728 : STD_LOGIC; 
  signal sig00000729 : STD_LOGIC; 
  signal sig0000072a : STD_LOGIC; 
  signal sig0000072b : STD_LOGIC; 
  signal sig0000072c : STD_LOGIC; 
  signal sig0000072d : STD_LOGIC; 
  signal sig0000072e : STD_LOGIC; 
  signal sig0000072f : STD_LOGIC; 
  signal sig00000730 : STD_LOGIC; 
  signal sig00000731 : STD_LOGIC; 
  signal sig00000732 : STD_LOGIC; 
  signal sig00000733 : STD_LOGIC; 
  signal sig00000734 : STD_LOGIC; 
  signal sig00000735 : STD_LOGIC; 
  signal sig00000736 : STD_LOGIC; 
  signal sig00000737 : STD_LOGIC; 
  signal sig00000738 : STD_LOGIC; 
  signal sig00000739 : STD_LOGIC; 
  signal sig0000073a : STD_LOGIC; 
  signal sig0000073b : STD_LOGIC; 
  signal sig0000073c : STD_LOGIC; 
  signal sig0000073d : STD_LOGIC; 
  signal sig0000073e : STD_LOGIC; 
  signal sig0000073f : STD_LOGIC; 
  signal sig00000740 : STD_LOGIC; 
  signal sig00000741 : STD_LOGIC; 
  signal sig00000742 : STD_LOGIC; 
  signal sig00000743 : STD_LOGIC; 
  signal sig00000744 : STD_LOGIC; 
  signal sig00000745 : STD_LOGIC; 
  signal sig00000746 : STD_LOGIC; 
  signal sig00000747 : STD_LOGIC; 
  signal sig00000748 : STD_LOGIC; 
  signal sig00000749 : STD_LOGIC; 
  signal sig0000074a : STD_LOGIC; 
  signal sig0000074b : STD_LOGIC; 
  signal sig0000074c : STD_LOGIC; 
  signal sig0000074d : STD_LOGIC; 
  signal sig0000074e : STD_LOGIC; 
  signal sig0000074f : STD_LOGIC; 
  signal sig00000750 : STD_LOGIC; 
  signal sig00000751 : STD_LOGIC; 
  signal sig00000752 : STD_LOGIC; 
  signal sig00000753 : STD_LOGIC; 
  signal sig00000754 : STD_LOGIC; 
  signal sig00000755 : STD_LOGIC; 
  signal sig00000756 : STD_LOGIC; 
  signal sig00000757 : STD_LOGIC; 
  signal sig00000758 : STD_LOGIC; 
  signal sig00000759 : STD_LOGIC; 
  signal sig0000075a : STD_LOGIC; 
  signal sig0000075b : STD_LOGIC; 
  signal sig0000075c : STD_LOGIC; 
  signal sig0000075d : STD_LOGIC; 
  signal sig0000075e : STD_LOGIC; 
  signal sig0000075f : STD_LOGIC; 
  signal sig00000760 : STD_LOGIC; 
  signal sig00000761 : STD_LOGIC; 
  signal sig00000762 : STD_LOGIC; 
  signal sig00000763 : STD_LOGIC; 
  signal sig00000764 : STD_LOGIC; 
  signal sig00000765 : STD_LOGIC; 
  signal sig00000766 : STD_LOGIC; 
  signal sig00000767 : STD_LOGIC; 
  signal sig00000768 : STD_LOGIC; 
  signal sig00000769 : STD_LOGIC; 
  signal sig0000076a : STD_LOGIC; 
  signal sig0000076b : STD_LOGIC; 
  signal sig0000076c : STD_LOGIC; 
  signal sig0000076d : STD_LOGIC; 
  signal sig0000076e : STD_LOGIC; 
  signal sig0000076f : STD_LOGIC; 
  signal sig00000770 : STD_LOGIC; 
  signal sig00000771 : STD_LOGIC; 
  signal sig00000772 : STD_LOGIC; 
  signal sig00000773 : STD_LOGIC; 
  signal sig00000774 : STD_LOGIC; 
  signal sig00000775 : STD_LOGIC; 
  signal sig00000776 : STD_LOGIC; 
  signal sig00000777 : STD_LOGIC; 
  signal sig00000778 : STD_LOGIC; 
  signal sig00000779 : STD_LOGIC; 
  signal sig0000077a : STD_LOGIC; 
  signal sig0000077b : STD_LOGIC; 
  signal sig0000077c : STD_LOGIC; 
  signal sig0000077d : STD_LOGIC; 
  signal sig0000077e : STD_LOGIC; 
  signal sig0000077f : STD_LOGIC; 
  signal sig00000780 : STD_LOGIC; 
  signal sig00000781 : STD_LOGIC; 
  signal sig00000782 : STD_LOGIC; 
  signal sig00000783 : STD_LOGIC; 
  signal sig00000784 : STD_LOGIC; 
  signal sig00000785 : STD_LOGIC; 
  signal sig00000786 : STD_LOGIC; 
  signal sig00000787 : STD_LOGIC; 
  signal sig00000788 : STD_LOGIC; 
  signal sig00000789 : STD_LOGIC; 
  signal sig0000078a : STD_LOGIC; 
  signal sig0000078b : STD_LOGIC; 
  signal sig0000078c : STD_LOGIC; 
  signal sig0000078d : STD_LOGIC; 
  signal sig0000078e : STD_LOGIC; 
  signal sig0000078f : STD_LOGIC; 
  signal sig00000790 : STD_LOGIC; 
  signal sig00000791 : STD_LOGIC; 
  signal sig00000792 : STD_LOGIC; 
  signal sig00000793 : STD_LOGIC; 
  signal sig00000794 : STD_LOGIC; 
  signal sig00000795 : STD_LOGIC; 
  signal sig00000796 : STD_LOGIC; 
  signal sig00000797 : STD_LOGIC; 
  signal sig00000798 : STD_LOGIC; 
  signal sig00000799 : STD_LOGIC; 
  signal sig0000079a : STD_LOGIC; 
  signal sig0000079b : STD_LOGIC; 
  signal sig0000079c : STD_LOGIC; 
  signal sig0000079d : STD_LOGIC; 
  signal sig0000079e : STD_LOGIC; 
  signal sig0000079f : STD_LOGIC; 
  signal sig000007a0 : STD_LOGIC; 
  signal sig000007a1 : STD_LOGIC; 
  signal sig000007a2 : STD_LOGIC; 
  signal sig000007a3 : STD_LOGIC; 
  signal sig000007a4 : STD_LOGIC; 
  signal sig000007a5 : STD_LOGIC; 
  signal sig000007a6 : STD_LOGIC; 
  signal sig000007a7 : STD_LOGIC; 
  signal sig000007a8 : STD_LOGIC; 
  signal sig000007a9 : STD_LOGIC; 
  signal sig000007aa : STD_LOGIC; 
  signal sig000007ab : STD_LOGIC; 
  signal sig000007ac : STD_LOGIC; 
  signal sig000007ad : STD_LOGIC; 
  signal sig000007ae : STD_LOGIC; 
  signal sig000007af : STD_LOGIC; 
  signal sig000007b0 : STD_LOGIC; 
  signal sig000007b1 : STD_LOGIC; 
  signal sig000007b2 : STD_LOGIC; 
  signal sig000007b3 : STD_LOGIC; 
  signal sig000007b4 : STD_LOGIC; 
  signal sig000007b5 : STD_LOGIC; 
  signal sig000007b6 : STD_LOGIC; 
  signal sig000007b7 : STD_LOGIC; 
  signal sig000007b8 : STD_LOGIC; 
  signal sig000007b9 : STD_LOGIC; 
  signal sig000007ba : STD_LOGIC; 
  signal sig000007bb : STD_LOGIC; 
  signal sig000007bc : STD_LOGIC; 
  signal sig000007bd : STD_LOGIC; 
  signal sig000007be : STD_LOGIC; 
  signal sig000007bf : STD_LOGIC; 
  signal sig000007c0 : STD_LOGIC; 
  signal sig000007c1 : STD_LOGIC; 
  signal sig000007c2 : STD_LOGIC; 
  signal sig000007c3 : STD_LOGIC; 
  signal sig000007c4 : STD_LOGIC; 
  signal sig000007c5 : STD_LOGIC; 
  signal sig000007c6 : STD_LOGIC; 
  signal sig000007c7 : STD_LOGIC; 
  signal sig000007c8 : STD_LOGIC; 
  signal sig000007c9 : STD_LOGIC; 
  signal sig000007ca : STD_LOGIC; 
  signal sig000007cb : STD_LOGIC; 
  signal sig000007cc : STD_LOGIC; 
  signal sig000007cd : STD_LOGIC; 
  signal sig000007ce : STD_LOGIC; 
  signal sig000007cf : STD_LOGIC; 
  signal sig000007d0 : STD_LOGIC; 
  signal sig000007d1 : STD_LOGIC; 
  signal sig000007d2 : STD_LOGIC; 
  signal sig000007d3 : STD_LOGIC; 
  signal sig000007d4 : STD_LOGIC; 
  signal sig000007d5 : STD_LOGIC; 
  signal sig000007d6 : STD_LOGIC; 
  signal sig000007d7 : STD_LOGIC; 
  signal sig000007d8 : STD_LOGIC; 
  signal sig000007d9 : STD_LOGIC; 
  signal sig000007da : STD_LOGIC; 
  signal sig000007db : STD_LOGIC; 
  signal sig000007dc : STD_LOGIC; 
  signal sig000007dd : STD_LOGIC; 
  signal sig000007de : STD_LOGIC; 
  signal sig000007df : STD_LOGIC; 
  signal sig000007e0 : STD_LOGIC; 
  signal sig000007e1 : STD_LOGIC; 
  signal sig000007e2 : STD_LOGIC; 
  signal sig000007e3 : STD_LOGIC; 
  signal sig000007e4 : STD_LOGIC; 
  signal sig000007e5 : STD_LOGIC; 
  signal sig000007e6 : STD_LOGIC; 
  signal sig000007e7 : STD_LOGIC; 
  signal sig000007e8 : STD_LOGIC; 
  signal sig000007e9 : STD_LOGIC; 
  signal sig000007ea : STD_LOGIC; 
  signal sig000007eb : STD_LOGIC; 
  signal sig000007ec : STD_LOGIC; 
  signal sig000007ed : STD_LOGIC; 
  signal sig000007ee : STD_LOGIC; 
  signal sig000007ef : STD_LOGIC; 
  signal sig000007f0 : STD_LOGIC; 
  signal sig000007f1 : STD_LOGIC; 
  signal sig000007f2 : STD_LOGIC; 
  signal sig000007f3 : STD_LOGIC; 
  signal sig000007f4 : STD_LOGIC; 
  signal sig000007f5 : STD_LOGIC; 
  signal sig000007f6 : STD_LOGIC; 
  signal sig000007f7 : STD_LOGIC; 
  signal sig000007f8 : STD_LOGIC; 
  signal sig000007f9 : STD_LOGIC; 
  signal sig000007fa : STD_LOGIC; 
  signal sig000007fb : STD_LOGIC; 
  signal sig000007fc : STD_LOGIC; 
  signal sig000007fd : STD_LOGIC; 
  signal sig000007fe : STD_LOGIC; 
  signal sig000007ff : STD_LOGIC; 
  signal sig00000800 : STD_LOGIC; 
  signal sig00000801 : STD_LOGIC; 
  signal sig00000802 : STD_LOGIC; 
  signal sig00000803 : STD_LOGIC; 
  signal sig00000804 : STD_LOGIC; 
  signal sig00000805 : STD_LOGIC; 
  signal sig00000806 : STD_LOGIC; 
  signal sig00000807 : STD_LOGIC; 
  signal sig00000808 : STD_LOGIC; 
  signal sig00000809 : STD_LOGIC; 
  signal sig0000080a : STD_LOGIC; 
  signal sig0000080b : STD_LOGIC; 
  signal sig0000080c : STD_LOGIC; 
  signal sig0000080d : STD_LOGIC; 
  signal sig0000080e : STD_LOGIC; 
  signal sig0000080f : STD_LOGIC; 
  signal sig00000810 : STD_LOGIC; 
  signal sig00000811 : STD_LOGIC; 
  signal sig00000812 : STD_LOGIC; 
  signal sig00000813 : STD_LOGIC; 
  signal sig00000814 : STD_LOGIC; 
  signal sig00000815 : STD_LOGIC; 
  signal sig00000816 : STD_LOGIC; 
  signal sig00000817 : STD_LOGIC; 
  signal sig00000818 : STD_LOGIC; 
  signal sig00000819 : STD_LOGIC; 
  signal sig0000081a : STD_LOGIC; 
  signal sig0000081b : STD_LOGIC; 
  signal sig0000081c : STD_LOGIC; 
  signal sig0000081d : STD_LOGIC; 
  signal sig0000081e : STD_LOGIC; 
  signal sig0000081f : STD_LOGIC; 
  signal sig00000820 : STD_LOGIC; 
  signal sig00000821 : STD_LOGIC; 
  signal sig00000822 : STD_LOGIC; 
  signal sig00000823 : STD_LOGIC; 
  signal sig00000824 : STD_LOGIC; 
  signal sig00000825 : STD_LOGIC; 
  signal sig00000826 : STD_LOGIC; 
  signal sig00000827 : STD_LOGIC; 
  signal sig00000828 : STD_LOGIC; 
  signal sig00000829 : STD_LOGIC; 
  signal sig0000082a : STD_LOGIC; 
  signal sig0000082b : STD_LOGIC; 
  signal sig0000082c : STD_LOGIC; 
  signal sig0000082d : STD_LOGIC; 
  signal sig0000082e : STD_LOGIC; 
  signal sig0000082f : STD_LOGIC; 
  signal sig00000830 : STD_LOGIC; 
  signal sig00000831 : STD_LOGIC; 
  signal sig00000832 : STD_LOGIC; 
  signal sig00000833 : STD_LOGIC; 
  signal sig00000834 : STD_LOGIC; 
  signal sig00000835 : STD_LOGIC; 
  signal sig00000836 : STD_LOGIC; 
  signal sig00000837 : STD_LOGIC; 
  signal sig00000838 : STD_LOGIC; 
  signal sig00000839 : STD_LOGIC; 
  signal sig0000083a : STD_LOGIC; 
  signal sig0000083b : STD_LOGIC; 
  signal sig0000083c : STD_LOGIC; 
  signal sig0000083d : STD_LOGIC; 
  signal sig0000083e : STD_LOGIC; 
  signal sig0000083f : STD_LOGIC; 
  signal sig00000840 : STD_LOGIC; 
  signal sig00000841 : STD_LOGIC; 
  signal sig00000842 : STD_LOGIC; 
  signal sig00000843 : STD_LOGIC; 
  signal sig00000844 : STD_LOGIC; 
  signal sig00000845 : STD_LOGIC; 
  signal sig00000846 : STD_LOGIC; 
  signal sig00000847 : STD_LOGIC; 
  signal sig00000848 : STD_LOGIC; 
  signal sig00000849 : STD_LOGIC; 
  signal sig0000084a : STD_LOGIC; 
  signal sig0000084b : STD_LOGIC; 
  signal sig0000084c : STD_LOGIC; 
  signal sig0000084d : STD_LOGIC; 
  signal sig0000084e : STD_LOGIC; 
  signal sig0000084f : STD_LOGIC; 
  signal sig00000850 : STD_LOGIC; 
  signal sig00000851 : STD_LOGIC; 
  signal sig00000852 : STD_LOGIC; 
  signal sig00000853 : STD_LOGIC; 
  signal sig00000854 : STD_LOGIC; 
  signal sig00000855 : STD_LOGIC; 
  signal sig00000856 : STD_LOGIC; 
  signal sig00000857 : STD_LOGIC; 
  signal sig00000858 : STD_LOGIC; 
  signal sig00000859 : STD_LOGIC; 
  signal sig0000085a : STD_LOGIC; 
  signal sig0000085b : STD_LOGIC; 
  signal sig0000085c : STD_LOGIC; 
  signal sig0000085d : STD_LOGIC; 
  signal sig0000085e : STD_LOGIC; 
  signal sig0000085f : STD_LOGIC; 
  signal sig00000860 : STD_LOGIC; 
  signal sig00000861 : STD_LOGIC; 
  signal sig00000862 : STD_LOGIC; 
  signal sig00000863 : STD_LOGIC; 
  signal sig00000864 : STD_LOGIC; 
  signal sig00000865 : STD_LOGIC; 
  signal sig00000866 : STD_LOGIC; 
  signal sig00000867 : STD_LOGIC; 
  signal sig00000868 : STD_LOGIC; 
  signal sig00000869 : STD_LOGIC; 
  signal sig0000086a : STD_LOGIC; 
  signal sig0000086b : STD_LOGIC; 
  signal sig0000086c : STD_LOGIC; 
  signal sig0000086d : STD_LOGIC; 
  signal sig0000086e : STD_LOGIC; 
  signal sig0000086f : STD_LOGIC; 
  signal sig00000870 : STD_LOGIC; 
  signal sig00000871 : STD_LOGIC; 
  signal sig00000872 : STD_LOGIC; 
  signal sig00000873 : STD_LOGIC; 
  signal sig00000874 : STD_LOGIC; 
  signal sig00000875 : STD_LOGIC; 
  signal sig00000876 : STD_LOGIC; 
  signal sig00000877 : STD_LOGIC; 
  signal sig00000878 : STD_LOGIC; 
  signal sig00000879 : STD_LOGIC; 
  signal sig0000087a : STD_LOGIC; 
  signal sig0000087b : STD_LOGIC; 
  signal sig0000087c : STD_LOGIC; 
  signal sig0000087d : STD_LOGIC; 
  signal sig0000087e : STD_LOGIC; 
  signal sig0000087f : STD_LOGIC; 
  signal sig00000880 : STD_LOGIC; 
  signal sig00000881 : STD_LOGIC; 
  signal sig00000882 : STD_LOGIC; 
  signal sig00000883 : STD_LOGIC; 
  signal sig00000884 : STD_LOGIC; 
  signal sig00000885 : STD_LOGIC; 
  signal sig00000886 : STD_LOGIC; 
  signal sig00000887 : STD_LOGIC; 
  signal sig00000888 : STD_LOGIC; 
  signal sig00000889 : STD_LOGIC; 
  signal sig0000088a : STD_LOGIC; 
  signal sig0000088b : STD_LOGIC; 
  signal sig0000088c : STD_LOGIC; 
  signal sig0000088d : STD_LOGIC; 
  signal sig0000088e : STD_LOGIC; 
  signal sig0000088f : STD_LOGIC; 
  signal sig00000890 : STD_LOGIC; 
  signal sig00000891 : STD_LOGIC; 
  signal sig00000892 : STD_LOGIC; 
  signal sig00000893 : STD_LOGIC; 
  signal sig00000894 : STD_LOGIC; 
  signal sig00000895 : STD_LOGIC; 
  signal sig00000896 : STD_LOGIC; 
  signal sig00000897 : STD_LOGIC; 
  signal sig00000898 : STD_LOGIC; 
  signal sig00000899 : STD_LOGIC; 
  signal sig0000089a : STD_LOGIC; 
  signal sig0000089b : STD_LOGIC; 
  signal sig0000089c : STD_LOGIC; 
  signal sig0000089d : STD_LOGIC; 
  signal sig0000089e : STD_LOGIC; 
  signal sig0000089f : STD_LOGIC; 
  signal sig000008a0 : STD_LOGIC; 
  signal sig000008a1 : STD_LOGIC; 
  signal sig000008a2 : STD_LOGIC; 
  signal sig000008a3 : STD_LOGIC; 
  signal sig000008b6 : STD_LOGIC; 
  signal sig000008cf : STD_LOGIC; 
  signal sig000008d0 : STD_LOGIC; 
  signal sig000008d1 : STD_LOGIC; 
  signal sig000008d2 : STD_LOGIC; 
  signal sig000008d3 : STD_LOGIC; 
  signal sig000008d4 : STD_LOGIC; 
  signal sig000008d5 : STD_LOGIC; 
  signal sig000008d6 : STD_LOGIC; 
  signal sig000008d7 : STD_LOGIC; 
  signal sig000008d8 : STD_LOGIC; 
  signal sig000008d9 : STD_LOGIC; 
  signal sig000008da : STD_LOGIC; 
  signal sig000008db : STD_LOGIC; 
  signal sig000008dc : STD_LOGIC; 
  signal sig000008dd : STD_LOGIC; 
  signal sig000008de : STD_LOGIC; 
  signal sig000008df : STD_LOGIC; 
  signal sig000008e0 : STD_LOGIC; 
  signal sig000008e1 : STD_LOGIC; 
  signal sig000008e2 : STD_LOGIC; 
  signal sig000008e3 : STD_LOGIC; 
  signal sig000008e4 : STD_LOGIC; 
  signal sig000008e5 : STD_LOGIC; 
  signal sig000008e6 : STD_LOGIC; 
  signal sig000008e7 : STD_LOGIC; 
  signal sig000008e8 : STD_LOGIC; 
  signal sig000008e9 : STD_LOGIC; 
  signal sig000008ea : STD_LOGIC; 
  signal sig000008eb : STD_LOGIC; 
  signal sig000008ec : STD_LOGIC; 
  signal sig000008ed : STD_LOGIC; 
  signal sig000008ee : STD_LOGIC; 
  signal sig000008ef : STD_LOGIC; 
  signal sig000008f0 : STD_LOGIC; 
  signal sig000008f1 : STD_LOGIC; 
  signal sig000008f2 : STD_LOGIC; 
  signal sig000008f3 : STD_LOGIC; 
  signal sig000008f4 : STD_LOGIC; 
  signal sig000008f5 : STD_LOGIC; 
  signal sig000008f6 : STD_LOGIC; 
  signal sig000008f7 : STD_LOGIC; 
  signal sig000008f8 : STD_LOGIC; 
  signal sig000008f9 : STD_LOGIC; 
  signal sig00000941 : STD_LOGIC; 
  signal sig00000942 : STD_LOGIC; 
  signal sig00000943 : STD_LOGIC; 
  signal sig00000944 : STD_LOGIC; 
  signal sig00000945 : STD_LOGIC; 
  signal sig00000946 : STD_LOGIC; 
  signal sig00000947 : STD_LOGIC; 
  signal sig00000948 : STD_LOGIC; 
  signal sig00000949 : STD_LOGIC; 
  signal sig0000094a : STD_LOGIC; 
  signal sig0000094b : STD_LOGIC; 
  signal sig0000094c : STD_LOGIC; 
  signal sig0000094d : STD_LOGIC; 
  signal sig0000094e : STD_LOGIC; 
  signal sig0000094f : STD_LOGIC; 
  signal sig0000097b : STD_LOGIC; 
  signal sig0000097c : STD_LOGIC; 
  signal sig0000097d : STD_LOGIC; 
  signal sig0000097e : STD_LOGIC; 
  signal sig0000097f : STD_LOGIC; 
  signal sig00000980 : STD_LOGIC; 
  signal sig00000981 : STD_LOGIC; 
  signal sig00000982 : STD_LOGIC; 
  signal sig00000983 : STD_LOGIC; 
  signal sig00000984 : STD_LOGIC; 
  signal sig00000985 : STD_LOGIC; 
  signal sig00000986 : STD_LOGIC; 
  signal sig00000987 : STD_LOGIC; 
  signal sig00000988 : STD_LOGIC; 
  signal sig00000989 : STD_LOGIC; 
  signal sig0000098a : STD_LOGIC; 
  signal sig0000098b : STD_LOGIC; 
  signal sig0000098c : STD_LOGIC; 
  signal sig0000098d : STD_LOGIC; 
  signal sig0000098e : STD_LOGIC; 
  signal sig0000098f : STD_LOGIC; 
  signal sig00000990 : STD_LOGIC; 
  signal sig00000991 : STD_LOGIC; 
  signal sig00000992 : STD_LOGIC; 
  signal sig00000993 : STD_LOGIC; 
  signal sig00000994 : STD_LOGIC; 
  signal sig00000995 : STD_LOGIC; 
  signal sig00000996 : STD_LOGIC; 
  signal sig00000997 : STD_LOGIC; 
  signal sig00000998 : STD_LOGIC; 
  signal sig00000999 : STD_LOGIC; 
  signal sig0000099a : STD_LOGIC; 
  signal sig0000099b : STD_LOGIC; 
  signal sig0000099c : STD_LOGIC; 
  signal sig0000099d : STD_LOGIC; 
  signal sig0000099e : STD_LOGIC; 
  signal sig0000099f : STD_LOGIC; 
  signal sig000009a0 : STD_LOGIC; 
  signal sig000009a1 : STD_LOGIC; 
  signal sig000009a2 : STD_LOGIC; 
  signal sig000009a3 : STD_LOGIC; 
  signal sig000009a4 : STD_LOGIC; 
  signal sig000009a5 : STD_LOGIC; 
  signal sig000009a7 : STD_LOGIC; 
  signal sig000009a8 : STD_LOGIC; 
  signal sig000009a9 : STD_LOGIC; 
  signal sig000009aa : STD_LOGIC; 
  signal sig000009ab : STD_LOGIC; 
  signal sig000009ac : STD_LOGIC; 
  signal sig000009ad : STD_LOGIC; 
  signal sig000009ae : STD_LOGIC; 
  signal sig000009af : STD_LOGIC; 
  signal sig000009b0 : STD_LOGIC; 
  signal sig000009b1 : STD_LOGIC; 
  signal sig000009b2 : STD_LOGIC; 
  signal sig000009b3 : STD_LOGIC; 
  signal sig000009b4 : STD_LOGIC; 
  signal sig000009b5 : STD_LOGIC; 
  signal sig000009b6 : STD_LOGIC; 
  signal sig000009b7 : STD_LOGIC; 
  signal sig000009b8 : STD_LOGIC; 
  signal sig000009b9 : STD_LOGIC; 
  signal sig000009ba : STD_LOGIC; 
  signal sig000009bb : STD_LOGIC; 
  signal sig000009bc : STD_LOGIC; 
  signal sig000009bd : STD_LOGIC; 
  signal sig000009be : STD_LOGIC; 
  signal sig000009bf : STD_LOGIC; 
  signal sig000009c0 : STD_LOGIC; 
  signal sig000009c1 : STD_LOGIC; 
  signal sig000009c2 : STD_LOGIC; 
  signal sig000009c3 : STD_LOGIC; 
  signal sig000009c4 : STD_LOGIC; 
  signal sig000009c5 : STD_LOGIC; 
  signal sig000009c6 : STD_LOGIC; 
  signal sig000009c7 : STD_LOGIC; 
  signal sig000009c8 : STD_LOGIC; 
  signal sig000009c9 : STD_LOGIC; 
  signal sig000009ca : STD_LOGIC; 
  signal sig000009cb : STD_LOGIC; 
  signal sig000009cc : STD_LOGIC; 
  signal sig000009cd : STD_LOGIC; 
  signal sig000009ce : STD_LOGIC; 
  signal sig000009cf : STD_LOGIC; 
  signal sig000009d0 : STD_LOGIC; 
  signal sig000009d1 : STD_LOGIC; 
  signal sig000009d2 : STD_LOGIC; 
  signal sig000009d3 : STD_LOGIC; 
  signal sig000009d4 : STD_LOGIC; 
  signal sig000009d5 : STD_LOGIC; 
  signal sig000009d6 : STD_LOGIC; 
  signal sig000009d7 : STD_LOGIC; 
  signal sig000009d8 : STD_LOGIC; 
  signal sig000009d9 : STD_LOGIC; 
  signal sig000009da : STD_LOGIC; 
  signal sig000009db : STD_LOGIC; 
  signal sig000009dc : STD_LOGIC; 
  signal sig000009dd : STD_LOGIC; 
  signal sig000009de : STD_LOGIC; 
  signal sig000009df : STD_LOGIC; 
  signal sig000009e0 : STD_LOGIC; 
  signal sig000009e1 : STD_LOGIC; 
  signal sig000009e2 : STD_LOGIC; 
  signal sig000009e3 : STD_LOGIC; 
  signal sig000009e4 : STD_LOGIC; 
  signal sig000009e5 : STD_LOGIC; 
  signal sig000009e6 : STD_LOGIC; 
  signal sig000009e7 : STD_LOGIC; 
  signal sig000009e8 : STD_LOGIC; 
  signal sig000009e9 : STD_LOGIC; 
  signal sig000009ea : STD_LOGIC; 
  signal sig000009eb : STD_LOGIC; 
  signal sig000009ec : STD_LOGIC; 
  signal sig000009ed : STD_LOGIC; 
  signal sig000009ee : STD_LOGIC; 
  signal sig000009ef : STD_LOGIC; 
  signal sig000009f0 : STD_LOGIC; 
  signal sig000009f1 : STD_LOGIC; 
  signal sig000009f2 : STD_LOGIC; 
  signal sig000009f3 : STD_LOGIC; 
  signal sig000009f4 : STD_LOGIC; 
  signal sig000009f5 : STD_LOGIC; 
  signal sig000009f6 : STD_LOGIC; 
  signal sig000009f7 : STD_LOGIC; 
  signal sig000009f8 : STD_LOGIC; 
  signal sig000009f9 : STD_LOGIC; 
  signal sig00000a22 : STD_LOGIC; 
  signal sig00000a23 : STD_LOGIC; 
  signal sig00000a24 : STD_LOGIC; 
  signal sig00000a25 : STD_LOGIC; 
  signal sig00000a28 : STD_LOGIC; 
  signal sig00000a29 : STD_LOGIC; 
  signal sig00000a2b : STD_LOGIC; 
  signal sig00000a2f : STD_LOGIC; 
  signal sig00000a35 : STD_LOGIC; 
  signal sig00000a36 : STD_LOGIC; 
  signal sig00000a37 : STD_LOGIC; 
  signal sig00000a38 : STD_LOGIC; 
  signal sig00000a39 : STD_LOGIC; 
  signal sig00000a3a : STD_LOGIC; 
  signal sig00000a3b : STD_LOGIC; 
  signal sig00000a3c : STD_LOGIC; 
  signal sig00000a3d : STD_LOGIC; 
  signal sig00000a3e : STD_LOGIC; 
  signal sig00000a3f : STD_LOGIC; 
  signal sig00000a40 : STD_LOGIC; 
  signal sig00000a41 : STD_LOGIC; 
  signal sig00000a42 : STD_LOGIC; 
  signal sig00000a43 : STD_LOGIC; 
  signal sig00000a44 : STD_LOGIC; 
  signal sig00000a45 : STD_LOGIC; 
  signal sig00000a46 : STD_LOGIC; 
  signal sig00000a47 : STD_LOGIC; 
  signal sig00000a48 : STD_LOGIC; 
  signal sig00000a49 : STD_LOGIC; 
  signal sig00000a4a : STD_LOGIC; 
  signal sig00000a4b : STD_LOGIC; 
  signal sig00000a4c : STD_LOGIC; 
  signal sig00000a4d : STD_LOGIC; 
  signal sig00000a4e : STD_LOGIC; 
  signal sig00000a4f : STD_LOGIC; 
  signal sig00000a50 : STD_LOGIC; 
  signal sig00000a51 : STD_LOGIC; 
  signal sig00000a52 : STD_LOGIC; 
  signal sig00000a53 : STD_LOGIC; 
  signal sig00000a54 : STD_LOGIC; 
  signal sig00000a55 : STD_LOGIC; 
  signal sig00000a56 : STD_LOGIC; 
  signal sig00000a57 : STD_LOGIC; 
  signal sig00000a58 : STD_LOGIC; 
  signal sig00000a59 : STD_LOGIC; 
  signal sig00000a5a : STD_LOGIC; 
  signal sig00000a5b : STD_LOGIC; 
  signal sig00000a5c : STD_LOGIC; 
  signal sig00000a5d : STD_LOGIC; 
  signal sig00000a5e : STD_LOGIC; 
  signal sig00000a5f : STD_LOGIC; 
  signal sig00000a60 : STD_LOGIC; 
  signal sig00000a61 : STD_LOGIC; 
  signal sig00000a62 : STD_LOGIC; 
  signal sig00000a63 : STD_LOGIC; 
  signal sig00000a64 : STD_LOGIC; 
  signal sig00000a65 : STD_LOGIC; 
  signal sig00000a66 : STD_LOGIC; 
  signal sig00000a67 : STD_LOGIC; 
  signal sig00000a68 : STD_LOGIC; 
  signal sig00000a69 : STD_LOGIC; 
  signal sig00000a6a : STD_LOGIC; 
  signal sig00000a6b : STD_LOGIC; 
  signal sig00000a6c : STD_LOGIC; 
  signal sig00000a6d : STD_LOGIC; 
  signal sig00000a6e : STD_LOGIC; 
  signal sig00000a6f : STD_LOGIC; 
  signal sig00000a70 : STD_LOGIC; 
  signal sig00000a71 : STD_LOGIC; 
  signal sig00000a72 : STD_LOGIC; 
  signal sig00000a73 : STD_LOGIC; 
  signal sig00000a74 : STD_LOGIC; 
  signal sig00000a75 : STD_LOGIC; 
  signal sig00000a76 : STD_LOGIC; 
  signal sig00000a77 : STD_LOGIC; 
  signal sig00000a78 : STD_LOGIC; 
  signal sig00000a79 : STD_LOGIC; 
  signal sig00000a7a : STD_LOGIC; 
  signal sig00000a7b : STD_LOGIC; 
  signal sig00000a7c : STD_LOGIC; 
  signal sig00000a7d : STD_LOGIC; 
  signal sig00000a7e : STD_LOGIC; 
  signal sig00000a7f : STD_LOGIC; 
  signal sig00000a80 : STD_LOGIC; 
  signal sig00000a81 : STD_LOGIC; 
  signal sig00000a82 : STD_LOGIC; 
  signal sig00000a83 : STD_LOGIC; 
  signal sig00000a84 : STD_LOGIC; 
  signal sig00000a85 : STD_LOGIC; 
  signal sig00000a86 : STD_LOGIC; 
  signal sig00000a87 : STD_LOGIC; 
  signal sig00000a88 : STD_LOGIC; 
  signal sig00000a89 : STD_LOGIC; 
  signal sig00000a8a : STD_LOGIC; 
  signal sig00000a8b : STD_LOGIC; 
  signal sig00000a8c : STD_LOGIC; 
  signal sig00000a8d : STD_LOGIC; 
  signal sig00000a8e : STD_LOGIC; 
  signal sig00000a8f : STD_LOGIC; 
  signal sig00000a90 : STD_LOGIC; 
  signal sig00000a91 : STD_LOGIC; 
  signal sig00000a92 : STD_LOGIC; 
  signal sig00000a93 : STD_LOGIC; 
  signal sig00000a94 : STD_LOGIC; 
  signal sig00000a95 : STD_LOGIC; 
  signal sig00000a96 : STD_LOGIC; 
  signal sig00000a97 : STD_LOGIC; 
  signal sig00000a98 : STD_LOGIC; 
  signal sig00000a99 : STD_LOGIC; 
  signal sig00000a9a : STD_LOGIC; 
  signal sig00000a9b : STD_LOGIC; 
  signal sig00000a9c : STD_LOGIC; 
  signal sig00000a9d : STD_LOGIC; 
  signal sig00000a9e : STD_LOGIC; 
  signal sig00000a9f : STD_LOGIC; 
  signal sig00000aa0 : STD_LOGIC; 
  signal sig00000aa1 : STD_LOGIC; 
  signal sig00000aa2 : STD_LOGIC; 
  signal sig00000aa3 : STD_LOGIC; 
  signal sig00000aa4 : STD_LOGIC; 
  signal sig00000aa5 : STD_LOGIC; 
  signal sig00000aa6 : STD_LOGIC; 
  signal sig00000aa7 : STD_LOGIC; 
  signal sig00000aa8 : STD_LOGIC; 
  signal sig00000aa9 : STD_LOGIC; 
  signal sig00000aaa : STD_LOGIC; 
  signal sig00000aab : STD_LOGIC; 
  signal sig00000aac : STD_LOGIC; 
  signal sig00000aad : STD_LOGIC; 
  signal sig00000aae : STD_LOGIC; 
  signal sig00000aaf : STD_LOGIC; 
  signal sig00000ab0 : STD_LOGIC; 
  signal sig00000ab1 : STD_LOGIC; 
  signal sig00000ab2 : STD_LOGIC; 
  signal sig00000ab3 : STD_LOGIC; 
  signal sig00000ab4 : STD_LOGIC; 
  signal sig00000ab5 : STD_LOGIC; 
  signal sig00000ab6 : STD_LOGIC; 
  signal sig00000ab7 : STD_LOGIC; 
  signal sig00000ab8 : STD_LOGIC; 
  signal sig00000ab9 : STD_LOGIC; 
  signal sig00000aba : STD_LOGIC; 
  signal sig00000abb : STD_LOGIC; 
  signal sig00000abc : STD_LOGIC; 
  signal sig00000abd : STD_LOGIC; 
  signal sig00000abe : STD_LOGIC; 
  signal sig00000abf : STD_LOGIC; 
  signal sig00000ac0 : STD_LOGIC; 
  signal sig00000ac1 : STD_LOGIC; 
  signal sig00000ac2 : STD_LOGIC; 
  signal sig00000ac3 : STD_LOGIC; 
  signal sig00000ac4 : STD_LOGIC; 
  signal sig00000ac5 : STD_LOGIC; 
  signal sig00000ac6 : STD_LOGIC; 
  signal sig00000ac7 : STD_LOGIC; 
  signal sig00000ac8 : STD_LOGIC; 
  signal sig00000ac9 : STD_LOGIC; 
  signal sig00000aca : STD_LOGIC; 
  signal sig00000acb : STD_LOGIC; 
  signal sig00000acc : STD_LOGIC; 
  signal sig00000acd : STD_LOGIC; 
  signal sig00000ace : STD_LOGIC; 
  signal sig00000acf : STD_LOGIC; 
  signal sig00000ad0 : STD_LOGIC; 
  signal sig00000ad1 : STD_LOGIC; 
  signal sig00000ad2 : STD_LOGIC; 
  signal sig00000ad3 : STD_LOGIC; 
  signal sig00000ad4 : STD_LOGIC; 
  signal sig00000ad5 : STD_LOGIC; 
  signal sig00000ad6 : STD_LOGIC; 
  signal sig00000ad7 : STD_LOGIC; 
  signal sig00000ad8 : STD_LOGIC; 
  signal sig00000ad9 : STD_LOGIC; 
  signal sig00000ada : STD_LOGIC; 
  signal sig00000adb : STD_LOGIC; 
  signal sig00000adc : STD_LOGIC; 
  signal sig00000add : STD_LOGIC; 
  signal sig00000ade : STD_LOGIC; 
  signal sig00000adf : STD_LOGIC; 
  signal sig00000ae0 : STD_LOGIC; 
  signal sig00000ae1 : STD_LOGIC; 
  signal sig00000ae2 : STD_LOGIC; 
  signal sig00000ae3 : STD_LOGIC; 
  signal sig00000ae4 : STD_LOGIC; 
  signal sig00000ae5 : STD_LOGIC; 
  signal sig00000ae6 : STD_LOGIC; 
  signal sig00000ae7 : STD_LOGIC; 
  signal sig00000ae8 : STD_LOGIC; 
  signal sig00000ae9 : STD_LOGIC; 
  signal sig00000aea : STD_LOGIC; 
  signal sig00000aeb : STD_LOGIC; 
  signal sig00000aec : STD_LOGIC; 
  signal sig00000aed : STD_LOGIC; 
  signal sig00000aee : STD_LOGIC; 
  signal sig00000aef : STD_LOGIC; 
  signal sig00000af0 : STD_LOGIC; 
  signal sig00000af1 : STD_LOGIC; 
  signal sig00000af2 : STD_LOGIC; 
  signal sig00000af3 : STD_LOGIC; 
  signal sig00000af4 : STD_LOGIC; 
  signal sig00000af5 : STD_LOGIC; 
  signal sig00000af6 : STD_LOGIC; 
  signal sig00000af7 : STD_LOGIC; 
  signal sig00000af8 : STD_LOGIC; 
  signal sig00000af9 : STD_LOGIC; 
  signal sig00000afa : STD_LOGIC; 
  signal sig00000afb : STD_LOGIC; 
  signal sig00000afc : STD_LOGIC; 
  signal sig00000afd : STD_LOGIC; 
  signal sig00000afe : STD_LOGIC; 
  signal sig00000aff : STD_LOGIC; 
  signal sig00000b00 : STD_LOGIC; 
  signal sig00000b01 : STD_LOGIC; 
  signal sig00000b02 : STD_LOGIC; 
  signal sig00000b03 : STD_LOGIC; 
  signal sig00000b04 : STD_LOGIC; 
  signal sig00000b05 : STD_LOGIC; 
  signal sig00000b06 : STD_LOGIC; 
  signal sig00000b07 : STD_LOGIC; 
  signal sig00000b08 : STD_LOGIC; 
  signal sig00000b09 : STD_LOGIC; 
  signal sig00000b0a : STD_LOGIC; 
  signal sig00000b0b : STD_LOGIC; 
  signal sig00000b0c : STD_LOGIC; 
  signal sig00000b0d : STD_LOGIC; 
  signal sig00000b0e : STD_LOGIC; 
  signal sig00000b0f : STD_LOGIC; 
  signal sig00000b10 : STD_LOGIC; 
  signal sig00000b11 : STD_LOGIC; 
  signal sig00000b12 : STD_LOGIC; 
  signal sig00000b13 : STD_LOGIC; 
  signal sig00000b14 : STD_LOGIC; 
  signal sig00000b15 : STD_LOGIC; 
  signal sig00000b16 : STD_LOGIC; 
  signal sig00000b17 : STD_LOGIC; 
  signal sig00000b18 : STD_LOGIC; 
  signal sig00000b19 : STD_LOGIC; 
  signal sig00000b1a : STD_LOGIC; 
  signal sig00000b1b : STD_LOGIC; 
  signal sig00000b1c : STD_LOGIC; 
  signal sig00000b1d : STD_LOGIC; 
  signal sig00000b1e : STD_LOGIC; 
  signal sig00000b1f : STD_LOGIC; 
  signal sig00000b20 : STD_LOGIC; 
  signal sig00000b21 : STD_LOGIC; 
  signal sig00000b22 : STD_LOGIC; 
  signal sig00000b23 : STD_LOGIC; 
  signal sig00000b24 : STD_LOGIC; 
  signal sig00000b25 : STD_LOGIC; 
  signal sig00000b26 : STD_LOGIC; 
  signal sig00000b27 : STD_LOGIC; 
  signal sig00000b28 : STD_LOGIC; 
  signal sig00000b29 : STD_LOGIC; 
  signal sig00000b2a : STD_LOGIC; 
  signal sig00000b2b : STD_LOGIC; 
  signal sig00000b2c : STD_LOGIC; 
  signal sig00000b2d : STD_LOGIC; 
  signal sig00000b2e : STD_LOGIC; 
  signal sig00000b2f : STD_LOGIC; 
  signal sig00000b30 : STD_LOGIC; 
  signal sig00000b31 : STD_LOGIC; 
  signal sig00000b32 : STD_LOGIC; 
  signal sig00000b33 : STD_LOGIC; 
  signal sig00000b34 : STD_LOGIC; 
  signal sig00000b35 : STD_LOGIC; 
  signal sig00000b36 : STD_LOGIC; 
  signal sig00000b37 : STD_LOGIC; 
  signal sig00000b38 : STD_LOGIC; 
  signal sig00000b39 : STD_LOGIC; 
  signal sig00000b3a : STD_LOGIC; 
  signal sig00000b3b : STD_LOGIC; 
  signal sig00000b3c : STD_LOGIC; 
  signal sig00000b3d : STD_LOGIC; 
  signal sig00000b3e : STD_LOGIC; 
  signal sig00000b3f : STD_LOGIC; 
  signal sig00000b40 : STD_LOGIC; 
  signal sig00000b41 : STD_LOGIC; 
  signal sig00000b42 : STD_LOGIC; 
  signal sig00000b43 : STD_LOGIC; 
  signal sig00000b44 : STD_LOGIC; 
  signal sig00000b45 : STD_LOGIC; 
  signal sig00000b46 : STD_LOGIC; 
  signal sig00000b47 : STD_LOGIC; 
  signal sig00000b48 : STD_LOGIC; 
  signal sig00000b49 : STD_LOGIC; 
  signal sig00000b4a : STD_LOGIC; 
  signal sig00000b4b : STD_LOGIC; 
  signal sig00000b4c : STD_LOGIC; 
  signal sig00000b4d : STD_LOGIC; 
  signal sig00000b4e : STD_LOGIC; 
  signal sig00000b4f : STD_LOGIC; 
  signal sig00000b50 : STD_LOGIC; 
  signal sig00000b51 : STD_LOGIC; 
  signal sig00000b52 : STD_LOGIC; 
  signal sig00000b53 : STD_LOGIC; 
  signal sig00000b54 : STD_LOGIC; 
  signal sig00000b55 : STD_LOGIC; 
  signal sig00000b56 : STD_LOGIC; 
  signal sig00000b57 : STD_LOGIC; 
  signal sig00000b58 : STD_LOGIC; 
  signal sig00000b59 : STD_LOGIC; 
  signal sig00000b5a : STD_LOGIC; 
  signal sig00000b5b : STD_LOGIC; 
  signal sig00000b5c : STD_LOGIC; 
  signal sig00000b5d : STD_LOGIC; 
  signal sig00000b5e : STD_LOGIC; 
  signal sig00000b5f : STD_LOGIC; 
  signal sig00000b60 : STD_LOGIC; 
  signal sig00000b61 : STD_LOGIC; 
  signal sig00000b62 : STD_LOGIC; 
  signal sig00000b63 : STD_LOGIC; 
  signal sig00000b64 : STD_LOGIC; 
  signal sig00000b65 : STD_LOGIC; 
  signal sig00000b66 : STD_LOGIC; 
  signal sig00000b67 : STD_LOGIC; 
  signal sig00000b68 : STD_LOGIC; 
  signal sig00000b69 : STD_LOGIC; 
  signal sig00000b6a : STD_LOGIC; 
  signal sig00000b6b : STD_LOGIC; 
  signal sig00000b6c : STD_LOGIC; 
  signal sig00000b6d : STD_LOGIC; 
  signal sig00000b6e : STD_LOGIC; 
  signal sig00000b6f : STD_LOGIC; 
  signal sig00000b70 : STD_LOGIC; 
  signal sig00000b71 : STD_LOGIC; 
  signal sig00000b72 : STD_LOGIC; 
  signal sig00000b73 : STD_LOGIC; 
  signal sig00000b74 : STD_LOGIC; 
  signal sig00000b75 : STD_LOGIC; 
  signal sig00000b76 : STD_LOGIC; 
  signal sig00000b77 : STD_LOGIC; 
  signal sig00000b78 : STD_LOGIC; 
  signal sig00000b79 : STD_LOGIC; 
  signal sig00000b7a : STD_LOGIC; 
  signal sig00000b7b : STD_LOGIC; 
  signal sig00000b7c : STD_LOGIC; 
  signal sig00000b7d : STD_LOGIC; 
  signal sig00000b7e : STD_LOGIC; 
  signal sig00000b7f : STD_LOGIC; 
  signal sig00000b80 : STD_LOGIC; 
  signal sig00000b81 : STD_LOGIC; 
  signal sig00000b82 : STD_LOGIC; 
  signal sig00000b83 : STD_LOGIC; 
  signal sig00000b84 : STD_LOGIC; 
  signal sig00000b85 : STD_LOGIC; 
  signal sig00000b86 : STD_LOGIC; 
  signal sig00000b87 : STD_LOGIC; 
  signal sig00000b88 : STD_LOGIC; 
  signal sig00000b89 : STD_LOGIC; 
  signal sig00000b8a : STD_LOGIC; 
  signal sig00000b8b : STD_LOGIC; 
  signal sig00000b8c : STD_LOGIC; 
  signal sig00000b8d : STD_LOGIC; 
  signal sig00000b8e : STD_LOGIC; 
  signal sig00000b8f : STD_LOGIC; 
  signal sig00000b90 : STD_LOGIC; 
  signal sig00000b91 : STD_LOGIC; 
  signal sig00000b92 : STD_LOGIC; 
  signal sig00000b93 : STD_LOGIC; 
  signal sig00000b94 : STD_LOGIC; 
  signal sig00000b95 : STD_LOGIC; 
  signal sig00000b96 : STD_LOGIC; 
  signal sig00000b97 : STD_LOGIC; 
  signal sig00000b98 : STD_LOGIC; 
  signal sig00000b99 : STD_LOGIC; 
  signal sig00000b9a : STD_LOGIC; 
  signal sig00000b9b : STD_LOGIC; 
  signal sig00000b9c : STD_LOGIC; 
  signal sig00000b9d : STD_LOGIC; 
  signal sig00000b9e : STD_LOGIC; 
  signal sig00000b9f : STD_LOGIC; 
  signal sig00000ba0 : STD_LOGIC; 
  signal sig00000ba1 : STD_LOGIC; 
  signal sig00000ba2 : STD_LOGIC; 
  signal sig00000ba3 : STD_LOGIC; 
  signal sig00000ba4 : STD_LOGIC; 
  signal sig00000ba5 : STD_LOGIC; 
  signal sig00000ba6 : STD_LOGIC; 
  signal sig00000ba7 : STD_LOGIC; 
  signal sig00000ba8 : STD_LOGIC; 
  signal sig00000ba9 : STD_LOGIC; 
  signal sig00000baa : STD_LOGIC; 
  signal sig00000bab : STD_LOGIC; 
  signal sig00000bac : STD_LOGIC; 
  signal sig00000bad : STD_LOGIC; 
  signal sig00000bae : STD_LOGIC; 
  signal sig00000baf : STD_LOGIC; 
  signal sig00000bb0 : STD_LOGIC; 
  signal sig00000bb1 : STD_LOGIC; 
  signal sig00000bb2 : STD_LOGIC; 
  signal sig00000bb3 : STD_LOGIC; 
  signal sig00000bb4 : STD_LOGIC; 
  signal sig00000bb5 : STD_LOGIC; 
  signal sig00000bb6 : STD_LOGIC; 
  signal sig00000bb7 : STD_LOGIC; 
  signal sig00000bb8 : STD_LOGIC; 
  signal sig00000bb9 : STD_LOGIC; 
  signal sig00000bba : STD_LOGIC; 
  signal sig00000bbb : STD_LOGIC; 
  signal sig00000bbc : STD_LOGIC; 
  signal sig00000bbd : STD_LOGIC; 
  signal sig00000bbe : STD_LOGIC; 
  signal sig00000bbf : STD_LOGIC; 
  signal sig00000bc0 : STD_LOGIC; 
  signal sig00000bc1 : STD_LOGIC; 
  signal sig00000bc2 : STD_LOGIC; 
  signal sig00000bc3 : STD_LOGIC; 
  signal sig00000bc4 : STD_LOGIC; 
  signal sig00000bc5 : STD_LOGIC; 
  signal sig00000bc6 : STD_LOGIC; 
  signal sig00000bc7 : STD_LOGIC; 
  signal sig00000bc8 : STD_LOGIC; 
  signal sig00000bc9 : STD_LOGIC; 
  signal sig00000bca : STD_LOGIC; 
  signal sig00000bcb : STD_LOGIC; 
  signal sig00000bcc : STD_LOGIC; 
  signal sig00000bcd : STD_LOGIC; 
  signal sig00000bce : STD_LOGIC; 
  signal sig00000bcf : STD_LOGIC; 
  signal sig00000bd0 : STD_LOGIC; 
  signal sig00000bd1 : STD_LOGIC; 
  signal sig00000bd2 : STD_LOGIC; 
  signal sig00000bd3 : STD_LOGIC; 
  signal sig00000bd4 : STD_LOGIC; 
  signal sig00000bd5 : STD_LOGIC; 
  signal sig00000bd6 : STD_LOGIC; 
  signal sig00000bd7 : STD_LOGIC; 
  signal sig00000bd8 : STD_LOGIC; 
  signal sig00000bd9 : STD_LOGIC; 
  signal sig00000bda : STD_LOGIC; 
  signal sig00000bdb : STD_LOGIC; 
  signal sig00000bdc : STD_LOGIC; 
  signal sig00000bdd : STD_LOGIC; 
  signal sig00000bde : STD_LOGIC; 
  signal sig00000bdf : STD_LOGIC; 
  signal sig00000be0 : STD_LOGIC; 
  signal sig00000be1 : STD_LOGIC; 
  signal sig00000be2 : STD_LOGIC; 
  signal sig00000be3 : STD_LOGIC; 
  signal sig00000be4 : STD_LOGIC; 
  signal sig00000be5 : STD_LOGIC; 
  signal sig00000be6 : STD_LOGIC; 
  signal sig00000be7 : STD_LOGIC; 
  signal sig00000be8 : STD_LOGIC; 
  signal sig00000be9 : STD_LOGIC; 
  signal sig00000bea : STD_LOGIC; 
  signal sig00000beb : STD_LOGIC; 
  signal sig00000bec : STD_LOGIC; 
  signal sig00000bed : STD_LOGIC; 
  signal sig00000bee : STD_LOGIC; 
  signal sig00000bef : STD_LOGIC; 
  signal sig00000bf0 : STD_LOGIC; 
  signal sig00000bf1 : STD_LOGIC; 
  signal sig00000bf2 : STD_LOGIC; 
  signal sig00000bf3 : STD_LOGIC; 
  signal sig00000bf4 : STD_LOGIC; 
  signal sig00000bf5 : STD_LOGIC; 
  signal sig00000bf6 : STD_LOGIC; 
  signal sig00000bf7 : STD_LOGIC; 
  signal sig00000bf8 : STD_LOGIC; 
  signal sig00000bf9 : STD_LOGIC; 
  signal sig00000bfa : STD_LOGIC; 
  signal sig00000bfb : STD_LOGIC; 
  signal sig00000bfc : STD_LOGIC; 
  signal sig00000bfd : STD_LOGIC; 
  signal sig00000bfe : STD_LOGIC; 
  signal sig00000bff : STD_LOGIC; 
  signal sig00000c00 : STD_LOGIC; 
  signal sig00000c01 : STD_LOGIC; 
  signal sig00000c02 : STD_LOGIC; 
  signal sig00000c03 : STD_LOGIC; 
  signal sig00000c04 : STD_LOGIC; 
  signal sig00000c05 : STD_LOGIC; 
  signal sig00000c06 : STD_LOGIC; 
  signal sig00000c07 : STD_LOGIC; 
  signal sig00000c08 : STD_LOGIC; 
  signal sig00000c09 : STD_LOGIC; 
  signal sig00000c0a : STD_LOGIC; 
  signal sig00000c0b : STD_LOGIC; 
  signal sig00000c0c : STD_LOGIC; 
  signal sig00000c0d : STD_LOGIC; 
  signal sig00000c0e : STD_LOGIC; 
  signal sig00000c0f : STD_LOGIC; 
  signal sig00000c10 : STD_LOGIC; 
  signal sig00000c11 : STD_LOGIC; 
  signal sig00000c12 : STD_LOGIC; 
  signal sig00000c13 : STD_LOGIC; 
  signal sig00000c14 : STD_LOGIC; 
  signal sig00000c15 : STD_LOGIC; 
  signal sig00000c16 : STD_LOGIC; 
  signal sig00000c17 : STD_LOGIC; 
  signal sig00000c18 : STD_LOGIC; 
  signal sig00000c19 : STD_LOGIC; 
  signal sig00000c1a : STD_LOGIC; 
  signal sig00000c1b : STD_LOGIC; 
  signal sig00000c1c : STD_LOGIC; 
  signal sig00000c1d : STD_LOGIC; 
  signal sig00000c1e : STD_LOGIC; 
  signal sig00000c1f : STD_LOGIC; 
  signal sig00000c20 : STD_LOGIC; 
  signal sig00000c21 : STD_LOGIC; 
  signal sig00000c22 : STD_LOGIC; 
  signal sig00000c23 : STD_LOGIC; 
  signal sig00000c24 : STD_LOGIC; 
  signal sig00000c25 : STD_LOGIC; 
  signal sig00000c26 : STD_LOGIC; 
  signal sig00000c27 : STD_LOGIC; 
  signal sig00000c28 : STD_LOGIC; 
  signal sig00000c29 : STD_LOGIC; 
  signal sig00000c2a : STD_LOGIC; 
  signal sig00000c2b : STD_LOGIC; 
  signal sig00000c2c : STD_LOGIC; 
  signal sig00000c2d : STD_LOGIC; 
  signal sig00000c2e : STD_LOGIC; 
  signal sig00000c2f : STD_LOGIC; 
  signal sig00000c30 : STD_LOGIC; 
  signal sig00000c31 : STD_LOGIC; 
  signal sig00000c32 : STD_LOGIC; 
  signal sig00000c33 : STD_LOGIC; 
  signal sig00000c34 : STD_LOGIC; 
  signal sig00000c35 : STD_LOGIC; 
  signal sig00000c36 : STD_LOGIC; 
  signal sig00000c37 : STD_LOGIC; 
  signal sig00000c38 : STD_LOGIC; 
  signal sig00000c39 : STD_LOGIC; 
  signal sig00000c3a : STD_LOGIC; 
  signal sig00000c3b : STD_LOGIC; 
  signal sig00000c3c : STD_LOGIC; 
  signal sig00000c3d : STD_LOGIC; 
  signal sig00000c3e : STD_LOGIC; 
  signal sig00000c3f : STD_LOGIC; 
  signal sig00000c40 : STD_LOGIC; 
  signal sig00000c41 : STD_LOGIC; 
  signal sig00000c42 : STD_LOGIC; 
  signal sig00000c43 : STD_LOGIC; 
  signal sig00000c44 : STD_LOGIC; 
  signal sig00000c45 : STD_LOGIC; 
  signal sig00000c46 : STD_LOGIC; 
  signal sig00000c47 : STD_LOGIC; 
  signal sig00000c48 : STD_LOGIC; 
  signal sig00000c49 : STD_LOGIC; 
  signal sig00000c4a : STD_LOGIC; 
  signal sig00000c4b : STD_LOGIC; 
  signal sig00000c4c : STD_LOGIC; 
  signal sig00000c4d : STD_LOGIC; 
  signal sig00000c4e : STD_LOGIC; 
  signal sig00000c4f : STD_LOGIC; 
  signal sig00000c50 : STD_LOGIC; 
  signal sig00000c51 : STD_LOGIC; 
  signal sig00000c52 : STD_LOGIC; 
  signal sig00000c53 : STD_LOGIC; 
  signal sig00000c54 : STD_LOGIC; 
  signal sig00000c55 : STD_LOGIC; 
  signal sig00000c56 : STD_LOGIC; 
  signal sig00000c57 : STD_LOGIC; 
  signal sig00000c58 : STD_LOGIC; 
  signal sig00000c59 : STD_LOGIC; 
  signal sig00000c5a : STD_LOGIC; 
  signal sig00000c5b : STD_LOGIC; 
  signal sig00000c5c : STD_LOGIC; 
  signal sig00000c5d : STD_LOGIC; 
  signal sig00000c5e : STD_LOGIC; 
  signal sig00000c5f : STD_LOGIC; 
  signal sig00000c60 : STD_LOGIC; 
  signal sig00000c61 : STD_LOGIC; 
  signal sig00000c62 : STD_LOGIC; 
  signal sig00000c63 : STD_LOGIC; 
  signal sig00000c64 : STD_LOGIC; 
  signal sig00000c65 : STD_LOGIC; 
  signal sig00000c66 : STD_LOGIC; 
  signal sig00000c67 : STD_LOGIC; 
  signal sig00000c68 : STD_LOGIC; 
  signal sig00000c69 : STD_LOGIC; 
  signal sig00000c6a : STD_LOGIC; 
  signal sig00000c6b : STD_LOGIC; 
  signal sig00000c6c : STD_LOGIC; 
  signal sig00000c6d : STD_LOGIC; 
  signal sig00000c6e : STD_LOGIC; 
  signal sig00000c6f : STD_LOGIC; 
  signal sig00000c70 : STD_LOGIC; 
  signal sig00000c71 : STD_LOGIC; 
  signal sig00000c72 : STD_LOGIC; 
  signal sig00000c73 : STD_LOGIC; 
  signal sig00000c74 : STD_LOGIC; 
  signal sig00000c75 : STD_LOGIC; 
  signal sig00000c76 : STD_LOGIC; 
  signal sig00000c77 : STD_LOGIC; 
  signal sig00000c78 : STD_LOGIC; 
  signal sig00000c79 : STD_LOGIC; 
  signal sig00000c7a : STD_LOGIC; 
  signal sig00000c7b : STD_LOGIC; 
  signal sig00000c7c : STD_LOGIC; 
  signal sig00000c7d : STD_LOGIC; 
  signal sig00000c7e : STD_LOGIC; 
  signal sig00000c7f : STD_LOGIC; 
  signal sig00000c80 : STD_LOGIC; 
  signal sig00000c81 : STD_LOGIC; 
  signal sig00000c82 : STD_LOGIC; 
  signal sig00000c83 : STD_LOGIC; 
  signal sig00000c84 : STD_LOGIC; 
  signal sig00000c85 : STD_LOGIC; 
  signal sig00000c86 : STD_LOGIC; 
  signal sig00000c87 : STD_LOGIC; 
  signal sig00000c88 : STD_LOGIC; 
  signal sig00000c89 : STD_LOGIC; 
  signal sig00000c8a : STD_LOGIC; 
  signal sig00000c8b : STD_LOGIC; 
  signal sig00000c8c : STD_LOGIC; 
  signal sig00000c8d : STD_LOGIC; 
  signal sig00000c8e : STD_LOGIC; 
  signal sig00000c8f : STD_LOGIC; 
  signal sig00000c90 : STD_LOGIC; 
  signal sig00000c91 : STD_LOGIC; 
  signal sig00000c92 : STD_LOGIC; 
  signal sig00000c93 : STD_LOGIC; 
  signal sig00000c94 : STD_LOGIC; 
  signal sig00000c95 : STD_LOGIC; 
  signal sig00000c96 : STD_LOGIC; 
  signal sig00000c97 : STD_LOGIC; 
  signal sig00000c98 : STD_LOGIC; 
  signal sig00000c99 : STD_LOGIC; 
  signal sig00000c9a : STD_LOGIC; 
  signal sig00000c9b : STD_LOGIC; 
  signal sig00000c9c : STD_LOGIC; 
  signal sig00000c9d : STD_LOGIC; 
  signal sig00000c9e : STD_LOGIC; 
  signal sig00000c9f : STD_LOGIC; 
  signal sig00000ca0 : STD_LOGIC; 
  signal sig00000ca1 : STD_LOGIC; 
  signal sig00000ca2 : STD_LOGIC; 
  signal sig00000ca3 : STD_LOGIC; 
  signal sig00000ca4 : STD_LOGIC; 
  signal sig00000ca5 : STD_LOGIC; 
  signal sig00000ca6 : STD_LOGIC; 
  signal sig00000ca7 : STD_LOGIC; 
  signal sig00000ca8 : STD_LOGIC; 
  signal sig00000ca9 : STD_LOGIC; 
  signal sig00000caa : STD_LOGIC; 
  signal sig00000cab : STD_LOGIC; 
  signal sig00000cac : STD_LOGIC; 
  signal sig00000cad : STD_LOGIC; 
  signal sig00000cae : STD_LOGIC; 
  signal sig00000caf : STD_LOGIC; 
  signal sig00000cb0 : STD_LOGIC; 
  signal sig00000cb1 : STD_LOGIC; 
  signal sig00000cb2 : STD_LOGIC; 
  signal sig00000cb3 : STD_LOGIC; 
  signal sig00000cb4 : STD_LOGIC; 
  signal sig00000cb5 : STD_LOGIC; 
  signal sig00000cb6 : STD_LOGIC; 
  signal sig00000cb7 : STD_LOGIC; 
  signal sig00000cb8 : STD_LOGIC; 
  signal sig00000cb9 : STD_LOGIC; 
  signal sig00000cba : STD_LOGIC; 
  signal sig00000cbb : STD_LOGIC; 
  signal sig00000cbc : STD_LOGIC; 
  signal sig00000cbd : STD_LOGIC; 
  signal sig00000cbe : STD_LOGIC; 
  signal sig00000cbf : STD_LOGIC; 
  signal sig00000cc0 : STD_LOGIC; 
  signal sig00000cc1 : STD_LOGIC; 
  signal sig00000cc2 : STD_LOGIC; 
  signal sig00000cc3 : STD_LOGIC; 
  signal sig00000cc4 : STD_LOGIC; 
  signal sig00000cc5 : STD_LOGIC; 
  signal sig00000cc6 : STD_LOGIC; 
  signal sig00000cc7 : STD_LOGIC; 
  signal sig00000cc8 : STD_LOGIC; 
  signal sig00000cc9 : STD_LOGIC; 
  signal sig00000cca : STD_LOGIC; 
  signal sig00000ccb : STD_LOGIC; 
  signal sig00000ccc : STD_LOGIC; 
  signal sig00000ccd : STD_LOGIC; 
  signal sig00000cce : STD_LOGIC; 
  signal sig00000ccf : STD_LOGIC; 
  signal sig00000cd0 : STD_LOGIC; 
  signal sig00000cd1 : STD_LOGIC; 
  signal sig00000cd2 : STD_LOGIC; 
  signal sig00000cd3 : STD_LOGIC; 
  signal sig00000cd4 : STD_LOGIC; 
  signal sig00000cd5 : STD_LOGIC; 
  signal sig00000cd6 : STD_LOGIC; 
  signal sig00000cd7 : STD_LOGIC; 
  signal sig00000cd8 : STD_LOGIC; 
  signal sig00000cd9 : STD_LOGIC; 
  signal sig00000cda : STD_LOGIC; 
  signal sig00000cdb : STD_LOGIC; 
  signal sig00000cdc : STD_LOGIC; 
  signal sig00000cdd : STD_LOGIC; 
  signal sig00000cde : STD_LOGIC; 
  signal sig00000cdf : STD_LOGIC; 
  signal sig00000ce0 : STD_LOGIC; 
  signal sig00000ce1 : STD_LOGIC; 
  signal sig00000ce2 : STD_LOGIC; 
  signal sig00000ce3 : STD_LOGIC; 
  signal sig00000ce4 : STD_LOGIC; 
  signal sig00000ce5 : STD_LOGIC; 
  signal sig00000ce6 : STD_LOGIC; 
  signal sig00000ce7 : STD_LOGIC; 
  signal sig00000ce8 : STD_LOGIC; 
  signal sig00000ce9 : STD_LOGIC; 
  signal sig00000cea : STD_LOGIC; 
  signal sig00000ceb : STD_LOGIC; 
  signal sig00000cec : STD_LOGIC; 
  signal sig00000ced : STD_LOGIC; 
  signal sig00000cee : STD_LOGIC; 
  signal sig00000cef : STD_LOGIC; 
  signal sig00000cf0 : STD_LOGIC; 
  signal sig00000cf1 : STD_LOGIC; 
  signal sig00000cf2 : STD_LOGIC; 
  signal sig00000cf3 : STD_LOGIC; 
  signal sig00000cf4 : STD_LOGIC; 
  signal sig00000cf5 : STD_LOGIC; 
  signal sig00000cf6 : STD_LOGIC; 
  signal sig00000cf7 : STD_LOGIC; 
  signal sig00000cf8 : STD_LOGIC; 
  signal sig00000cf9 : STD_LOGIC; 
  signal sig00000cfa : STD_LOGIC; 
  signal sig00000cfb : STD_LOGIC; 
  signal sig00000cfc : STD_LOGIC; 
  signal sig00000cfd : STD_LOGIC; 
  signal sig00000cfe : STD_LOGIC; 
  signal sig00000cff : STD_LOGIC; 
  signal sig00000d00 : STD_LOGIC; 
  signal sig00000d01 : STD_LOGIC; 
  signal sig00000d02 : STD_LOGIC; 
  signal sig00000d03 : STD_LOGIC; 
  signal sig00000d04 : STD_LOGIC; 
  signal sig00000d05 : STD_LOGIC; 
  signal sig00000d06 : STD_LOGIC; 
  signal sig00000d07 : STD_LOGIC; 
  signal sig00000d08 : STD_LOGIC; 
  signal sig00000d09 : STD_LOGIC; 
  signal sig00000d0a : STD_LOGIC; 
  signal sig00000d0b : STD_LOGIC; 
  signal sig00000d0c : STD_LOGIC; 
  signal sig00000d0d : STD_LOGIC; 
  signal sig00000d0e : STD_LOGIC; 
  signal sig00000d0f : STD_LOGIC; 
  signal sig00000d10 : STD_LOGIC; 
  signal sig00000d11 : STD_LOGIC; 
  signal sig00000d12 : STD_LOGIC; 
  signal sig00000d13 : STD_LOGIC; 
  signal sig00000d14 : STD_LOGIC; 
  signal sig00000d15 : STD_LOGIC; 
  signal sig00000d16 : STD_LOGIC; 
  signal sig00000d17 : STD_LOGIC; 
  signal sig00000d18 : STD_LOGIC; 
  signal sig00000d19 : STD_LOGIC; 
  signal sig00000d1a : STD_LOGIC; 
  signal sig00000d1b : STD_LOGIC; 
  signal sig00000d1c : STD_LOGIC; 
  signal sig00000d1d : STD_LOGIC; 
  signal sig00000d1e : STD_LOGIC; 
  signal sig00000d1f : STD_LOGIC; 
  signal sig00000d20 : STD_LOGIC; 
  signal sig00000d21 : STD_LOGIC; 
  signal sig00000d22 : STD_LOGIC; 
  signal sig00000d23 : STD_LOGIC; 
  signal sig00000d24 : STD_LOGIC; 
  signal sig00000d25 : STD_LOGIC; 
  signal sig00000d26 : STD_LOGIC; 
  signal sig00000d27 : STD_LOGIC; 
  signal sig00000d28 : STD_LOGIC; 
  signal sig00000d29 : STD_LOGIC; 
  signal sig00000d2a : STD_LOGIC; 
  signal sig00000d2b : STD_LOGIC; 
  signal sig00000d2c : STD_LOGIC; 
  signal sig00000d2d : STD_LOGIC; 
  signal sig00000d2e : STD_LOGIC; 
  signal sig00000d2f : STD_LOGIC; 
  signal sig00000d30 : STD_LOGIC; 
  signal sig00000d31 : STD_LOGIC; 
  signal sig00000d32 : STD_LOGIC; 
  signal sig00000d33 : STD_LOGIC; 
  signal sig00000d34 : STD_LOGIC; 
  signal sig00000d35 : STD_LOGIC; 
  signal sig00000d36 : STD_LOGIC; 
  signal sig00000d37 : STD_LOGIC; 
  signal sig00000d38 : STD_LOGIC; 
  signal sig00000d39 : STD_LOGIC; 
  signal sig00000d3a : STD_LOGIC; 
  signal sig00000d3b : STD_LOGIC; 
  signal sig00000d3c : STD_LOGIC; 
  signal sig00000d3d : STD_LOGIC; 
  signal sig00000d3e : STD_LOGIC; 
  signal sig00000d3f : STD_LOGIC; 
  signal sig00000d40 : STD_LOGIC; 
  signal sig00000d41 : STD_LOGIC; 
  signal sig00000d42 : STD_LOGIC; 
  signal sig00000d43 : STD_LOGIC; 
  signal sig00000d44 : STD_LOGIC; 
  signal sig00000d45 : STD_LOGIC; 
  signal sig00000d46 : STD_LOGIC; 
  signal sig00000d47 : STD_LOGIC; 
  signal sig00000d48 : STD_LOGIC; 
  signal sig00000d49 : STD_LOGIC; 
  signal sig00000d4a : STD_LOGIC; 
  signal sig00000d4b : STD_LOGIC; 
  signal sig00000d4c : STD_LOGIC; 
  signal sig00000d4d : STD_LOGIC; 
  signal sig00000d4e : STD_LOGIC; 
  signal sig00000d4f : STD_LOGIC; 
  signal sig00000d50 : STD_LOGIC; 
  signal sig00000d51 : STD_LOGIC; 
  signal sig00000d52 : STD_LOGIC; 
  signal sig00000d53 : STD_LOGIC; 
  signal sig00000d54 : STD_LOGIC; 
  signal sig00000d55 : STD_LOGIC; 
  signal sig00000d56 : STD_LOGIC; 
  signal sig00000d57 : STD_LOGIC; 
  signal sig00000d58 : STD_LOGIC; 
  signal sig00000d59 : STD_LOGIC; 
  signal sig00000d5a : STD_LOGIC; 
  signal sig00000d5b : STD_LOGIC; 
  signal sig00000d5c : STD_LOGIC; 
  signal sig00000d5d : STD_LOGIC; 
  signal sig00000d5e : STD_LOGIC; 
  signal sig00000d5f : STD_LOGIC; 
  signal sig00000d60 : STD_LOGIC; 
  signal sig00000d61 : STD_LOGIC; 
  signal sig00000d62 : STD_LOGIC; 
  signal sig00000d63 : STD_LOGIC; 
  signal sig00000d64 : STD_LOGIC; 
  signal sig00000d65 : STD_LOGIC; 
  signal sig00000d66 : STD_LOGIC; 
  signal sig00000d67 : STD_LOGIC; 
  signal sig00000d68 : STD_LOGIC; 
  signal sig00000d69 : STD_LOGIC; 
  signal sig00000d6a : STD_LOGIC; 
  signal sig00000d6b : STD_LOGIC; 
  signal sig00000d6c : STD_LOGIC; 
  signal sig00000d6d : STD_LOGIC; 
  signal sig00000d6e : STD_LOGIC; 
  signal sig00000d6f : STD_LOGIC; 
  signal sig00000d70 : STD_LOGIC; 
  signal sig00000d71 : STD_LOGIC; 
  signal sig00000d72 : STD_LOGIC; 
  signal sig00000d73 : STD_LOGIC; 
  signal sig00000d74 : STD_LOGIC; 
  signal sig00000d75 : STD_LOGIC; 
  signal sig00000d76 : STD_LOGIC; 
  signal sig00000d77 : STD_LOGIC; 
  signal sig00000d78 : STD_LOGIC; 
  signal sig00000d79 : STD_LOGIC; 
  signal sig00000d7a : STD_LOGIC; 
  signal sig00000d7b : STD_LOGIC; 
  signal sig00000d7c : STD_LOGIC; 
  signal sig00000d7d : STD_LOGIC; 
  signal sig00000d7e : STD_LOGIC; 
  signal sig00000d7f : STD_LOGIC; 
  signal sig00000d80 : STD_LOGIC; 
  signal sig00000d81 : STD_LOGIC; 
  signal sig00000d82 : STD_LOGIC; 
  signal sig00000d83 : STD_LOGIC; 
  signal sig00000d84 : STD_LOGIC; 
  signal sig00000d85 : STD_LOGIC; 
  signal sig00000d86 : STD_LOGIC; 
  signal sig00000d87 : STD_LOGIC; 
  signal sig00000d88 : STD_LOGIC; 
  signal sig00000d89 : STD_LOGIC; 
  signal sig00000d8a : STD_LOGIC; 
  signal sig00000d8b : STD_LOGIC; 
  signal sig00000d8c : STD_LOGIC; 
  signal sig00000d8d : STD_LOGIC; 
  signal sig00000d8e : STD_LOGIC; 
  signal sig00000d8f : STD_LOGIC; 
  signal sig00000d90 : STD_LOGIC; 
  signal sig00000d91 : STD_LOGIC; 
  signal sig00000d92 : STD_LOGIC; 
  signal sig00000d93 : STD_LOGIC; 
  signal sig00000d94 : STD_LOGIC; 
  signal sig00000d95 : STD_LOGIC; 
  signal sig00000d96 : STD_LOGIC; 
  signal sig00000d97 : STD_LOGIC; 
  signal sig00000d98 : STD_LOGIC; 
  signal sig00000d99 : STD_LOGIC; 
  signal sig00000d9a : STD_LOGIC; 
  signal sig00000d9b : STD_LOGIC; 
  signal sig00000d9c : STD_LOGIC; 
  signal sig00000d9d : STD_LOGIC; 
  signal sig00000d9e : STD_LOGIC; 
  signal sig00000d9f : STD_LOGIC; 
  signal sig00000da0 : STD_LOGIC; 
  signal sig00000da1 : STD_LOGIC; 
  signal sig00000da2 : STD_LOGIC; 
  signal sig00000da3 : STD_LOGIC; 
  signal sig00000da4 : STD_LOGIC; 
  signal sig00000da5 : STD_LOGIC; 
  signal sig00000da6 : STD_LOGIC; 
  signal sig00000da7 : STD_LOGIC; 
  signal sig00000da8 : STD_LOGIC; 
  signal sig00000da9 : STD_LOGIC; 
  signal sig00000daa : STD_LOGIC; 
  signal sig00000dab : STD_LOGIC; 
  signal sig00000dac : STD_LOGIC; 
  signal sig00000dad : STD_LOGIC; 
  signal sig00000dae : STD_LOGIC; 
  signal sig00000daf : STD_LOGIC; 
  signal sig00000db0 : STD_LOGIC; 
  signal sig00000db1 : STD_LOGIC; 
  signal sig00000db2 : STD_LOGIC; 
  signal sig00000db3 : STD_LOGIC; 
  signal sig00000db4 : STD_LOGIC; 
  signal sig00000db5 : STD_LOGIC; 
  signal sig00000db6 : STD_LOGIC; 
  signal sig00000db7 : STD_LOGIC; 
  signal sig00000db8 : STD_LOGIC; 
  signal sig00000db9 : STD_LOGIC; 
  signal sig00000dba : STD_LOGIC; 
  signal sig00000dbb : STD_LOGIC; 
  signal sig00000dbc : STD_LOGIC; 
  signal sig00000dbd : STD_LOGIC; 
  signal sig00000dbe : STD_LOGIC; 
  signal sig00000dbf : STD_LOGIC; 
  signal sig00000dc0 : STD_LOGIC; 
  signal sig00000dc1 : STD_LOGIC; 
  signal sig00000dc2 : STD_LOGIC; 
  signal sig00000dc3 : STD_LOGIC; 
  signal sig00000dc4 : STD_LOGIC; 
  signal sig00000dc5 : STD_LOGIC; 
  signal sig00000dc6 : STD_LOGIC; 
  signal sig00000dc7 : STD_LOGIC; 
  signal sig00000dc8 : STD_LOGIC; 
  signal sig00000dc9 : STD_LOGIC; 
  signal sig00000dca : STD_LOGIC; 
  signal sig00000dcb : STD_LOGIC; 
  signal sig00000dcc : STD_LOGIC; 
  signal sig00000dcd : STD_LOGIC; 
  signal sig00000dce : STD_LOGIC; 
  signal sig00000dcf : STD_LOGIC; 
  signal sig00000dd0 : STD_LOGIC; 
  signal sig00000dd1 : STD_LOGIC; 
  signal sig00000dd2 : STD_LOGIC; 
  signal sig00000dd3 : STD_LOGIC; 
  signal sig00000dd4 : STD_LOGIC; 
  signal sig00000dd5 : STD_LOGIC; 
  signal sig00000dd6 : STD_LOGIC; 
  signal sig00000dd7 : STD_LOGIC; 
  signal sig00000dd8 : STD_LOGIC; 
  signal sig00000dd9 : STD_LOGIC; 
  signal sig00000dda : STD_LOGIC; 
  signal sig00000ddb : STD_LOGIC; 
  signal sig00000ddc : STD_LOGIC; 
  signal sig00000ddd : STD_LOGIC; 
  signal sig00000dde : STD_LOGIC; 
  signal sig00000ddf : STD_LOGIC; 
  signal sig00000de0 : STD_LOGIC; 
  signal sig00000de1 : STD_LOGIC; 
  signal sig00000de2 : STD_LOGIC; 
  signal sig00000de3 : STD_LOGIC; 
  signal sig00000de4 : STD_LOGIC; 
  signal sig00000de5 : STD_LOGIC; 
  signal sig00000de6 : STD_LOGIC; 
  signal sig00000de7 : STD_LOGIC; 
  signal sig00000de8 : STD_LOGIC; 
  signal sig00000de9 : STD_LOGIC; 
  signal sig00000dea : STD_LOGIC; 
  signal sig00000deb : STD_LOGIC; 
  signal sig00000dec : STD_LOGIC; 
  signal sig00000ded : STD_LOGIC; 
  signal sig00000dee : STD_LOGIC; 
  signal sig00000def : STD_LOGIC; 
  signal sig00000df0 : STD_LOGIC; 
  signal sig00000df1 : STD_LOGIC; 
  signal sig00000df2 : STD_LOGIC; 
  signal sig00000df3 : STD_LOGIC; 
  signal sig00000df4 : STD_LOGIC; 
  signal sig00000df5 : STD_LOGIC; 
  signal sig00000df6 : STD_LOGIC; 
  signal sig00000df7 : STD_LOGIC; 
  signal sig00000df8 : STD_LOGIC; 
  signal sig00000df9 : STD_LOGIC; 
  signal sig00000dfa : STD_LOGIC; 
  signal sig00000dfb : STD_LOGIC; 
  signal sig00000dfc : STD_LOGIC; 
  signal sig00000dfd : STD_LOGIC; 
  signal sig00000dfe : STD_LOGIC; 
  signal sig00000dff : STD_LOGIC; 
  signal sig00000e00 : STD_LOGIC; 
  signal sig00000e01 : STD_LOGIC; 
  signal sig00000e02 : STD_LOGIC; 
  signal sig00000e03 : STD_LOGIC; 
  signal sig00000e04 : STD_LOGIC; 
  signal sig00000e05 : STD_LOGIC; 
  signal sig00000e06 : STD_LOGIC; 
  signal sig00000e07 : STD_LOGIC; 
  signal sig00000e08 : STD_LOGIC; 
  signal sig00000e09 : STD_LOGIC; 
  signal sig00000e0a : STD_LOGIC; 
  signal sig00000e0b : STD_LOGIC; 
  signal sig00000e0c : STD_LOGIC; 
  signal sig00000e0d : STD_LOGIC; 
  signal sig00000e0e : STD_LOGIC; 
  signal sig00000e0f : STD_LOGIC; 
  signal sig00000e10 : STD_LOGIC; 
  signal sig00000e11 : STD_LOGIC; 
  signal sig00000e12 : STD_LOGIC; 
  signal sig00000e13 : STD_LOGIC; 
  signal sig00000e14 : STD_LOGIC; 
  signal sig00000e15 : STD_LOGIC; 
  signal sig00000e16 : STD_LOGIC; 
  signal sig00000e17 : STD_LOGIC; 
  signal sig00000e18 : STD_LOGIC; 
  signal sig00000e19 : STD_LOGIC; 
  signal sig00000e1a : STD_LOGIC; 
  signal sig00000e1b : STD_LOGIC; 
  signal sig00000e1c : STD_LOGIC; 
  signal sig00000e1d : STD_LOGIC; 
  signal sig00000e1e : STD_LOGIC; 
  signal sig00000e1f : STD_LOGIC; 
  signal sig00000e20 : STD_LOGIC; 
  signal sig00000e21 : STD_LOGIC; 
  signal sig00000e22 : STD_LOGIC; 
  signal sig00000e23 : STD_LOGIC; 
  signal sig00000e24 : STD_LOGIC; 
  signal sig00000e25 : STD_LOGIC; 
  signal sig00000e26 : STD_LOGIC; 
  signal sig00000e27 : STD_LOGIC; 
  signal sig00000e28 : STD_LOGIC; 
  signal sig00000e29 : STD_LOGIC; 
  signal sig00000e2a : STD_LOGIC; 
  signal sig00000e2b : STD_LOGIC; 
  signal sig00000e2c : STD_LOGIC; 
  signal sig00000e2d : STD_LOGIC; 
  signal sig00000e2e : STD_LOGIC; 
  signal sig00000e2f : STD_LOGIC; 
  signal sig00000e30 : STD_LOGIC; 
  signal sig00000e31 : STD_LOGIC; 
  signal sig00000e32 : STD_LOGIC; 
  signal sig00000e33 : STD_LOGIC; 
  signal sig00000e34 : STD_LOGIC; 
  signal sig00000e35 : STD_LOGIC; 
  signal sig00000e36 : STD_LOGIC; 
  signal sig00000e37 : STD_LOGIC; 
  signal sig00000e38 : STD_LOGIC; 
  signal sig00000e39 : STD_LOGIC; 
  signal sig00000e3a : STD_LOGIC; 
  signal sig00000e3b : STD_LOGIC; 
  signal sig00000e3c : STD_LOGIC; 
  signal sig00000e3d : STD_LOGIC; 
  signal sig00000e3e : STD_LOGIC; 
  signal sig00000e3f : STD_LOGIC; 
  signal sig00000e40 : STD_LOGIC; 
  signal sig00000e41 : STD_LOGIC; 
  signal sig00000e42 : STD_LOGIC; 
  signal sig00000e43 : STD_LOGIC; 
  signal sig00000e44 : STD_LOGIC; 
  signal sig00000e45 : STD_LOGIC; 
  signal sig00000e46 : STD_LOGIC; 
  signal sig00000e47 : STD_LOGIC; 
  signal sig00000e48 : STD_LOGIC; 
  signal sig00000e49 : STD_LOGIC; 
  signal sig00000e4a : STD_LOGIC; 
  signal sig00000e4b : STD_LOGIC; 
  signal sig00000e4c : STD_LOGIC; 
  signal sig00000e4d : STD_LOGIC; 
  signal sig00000e4e : STD_LOGIC; 
  signal sig00000e4f : STD_LOGIC; 
  signal sig00000e50 : STD_LOGIC; 
  signal sig00000e51 : STD_LOGIC; 
  signal sig00000e52 : STD_LOGIC; 
  signal sig00000e53 : STD_LOGIC; 
  signal sig00000e54 : STD_LOGIC; 
  signal sig00000e55 : STD_LOGIC; 
  signal sig00000e56 : STD_LOGIC; 
  signal sig00000e57 : STD_LOGIC; 
  signal sig00000e58 : STD_LOGIC; 
  signal sig00000e59 : STD_LOGIC; 
  signal sig00000e5a : STD_LOGIC; 
  signal sig00000e5b : STD_LOGIC; 
  signal sig00000e5c : STD_LOGIC; 
  signal sig00000e5d : STD_LOGIC; 
  signal sig00000e5e : STD_LOGIC; 
  signal sig00000e5f : STD_LOGIC; 
  signal sig00000e60 : STD_LOGIC; 
  signal sig00000e61 : STD_LOGIC; 
  signal sig00000e62 : STD_LOGIC; 
  signal sig00000e63 : STD_LOGIC; 
  signal sig00000e64 : STD_LOGIC; 
  signal sig00000e65 : STD_LOGIC; 
  signal sig00000e66 : STD_LOGIC; 
  signal sig00000e67 : STD_LOGIC; 
  signal sig00000e68 : STD_LOGIC; 
  signal sig00000e69 : STD_LOGIC; 
  signal sig00000e6a : STD_LOGIC; 
  signal sig00000e6b : STD_LOGIC; 
  signal sig00000e6c : STD_LOGIC; 
  signal sig00000e6d : STD_LOGIC; 
  signal sig00000e6e : STD_LOGIC; 
  signal sig00000e6f : STD_LOGIC; 
  signal sig00000e70 : STD_LOGIC; 
  signal sig00000e71 : STD_LOGIC; 
  signal sig00000e72 : STD_LOGIC; 
  signal sig00000e73 : STD_LOGIC; 
  signal sig00000e74 : STD_LOGIC; 
  signal sig00000e75 : STD_LOGIC; 
  signal sig00000e76 : STD_LOGIC; 
  signal sig00000e77 : STD_LOGIC; 
  signal sig00000e78 : STD_LOGIC; 
  signal sig00000e79 : STD_LOGIC; 
  signal sig00000e7a : STD_LOGIC; 
  signal sig00000e7b : STD_LOGIC; 
  signal sig00000e7c : STD_LOGIC; 
  signal sig00000e7d : STD_LOGIC; 
  signal sig00000e7e : STD_LOGIC; 
  signal sig00000e7f : STD_LOGIC; 
  signal sig00000e80 : STD_LOGIC; 
  signal sig00000e81 : STD_LOGIC; 
  signal sig00000e82 : STD_LOGIC; 
  signal sig00000e83 : STD_LOGIC; 
  signal sig00000e84 : STD_LOGIC; 
  signal sig00000e85 : STD_LOGIC; 
  signal sig00000e86 : STD_LOGIC; 
  signal sig00000e87 : STD_LOGIC; 
  signal sig00000e88 : STD_LOGIC; 
  signal sig00000e89 : STD_LOGIC; 
  signal sig00000e8a : STD_LOGIC; 
  signal sig00000e8b : STD_LOGIC; 
  signal sig00000e8c : STD_LOGIC; 
  signal sig00000e8d : STD_LOGIC; 
  signal sig00000e8e : STD_LOGIC; 
  signal sig00000e8f : STD_LOGIC; 
  signal sig00000e90 : STD_LOGIC; 
  signal sig00000e91 : STD_LOGIC; 
  signal sig00000e92 : STD_LOGIC; 
  signal sig00000e93 : STD_LOGIC; 
  signal sig00000e94 : STD_LOGIC; 
  signal sig00000e95 : STD_LOGIC; 
  signal sig00000e96 : STD_LOGIC; 
  signal sig00000e97 : STD_LOGIC; 
  signal sig00000e98 : STD_LOGIC; 
  signal sig00000e99 : STD_LOGIC; 
  signal sig00000e9a : STD_LOGIC; 
  signal sig00000e9b : STD_LOGIC; 
  signal sig00000e9c : STD_LOGIC; 
  signal sig00000e9d : STD_LOGIC; 
  signal sig00000e9e : STD_LOGIC; 
  signal sig00000e9f : STD_LOGIC; 
  signal sig00000ea0 : STD_LOGIC; 
  signal sig00000ea1 : STD_LOGIC; 
  signal sig00000ea2 : STD_LOGIC; 
  signal sig00000ea3 : STD_LOGIC; 
  signal sig00000ea4 : STD_LOGIC; 
  signal sig00000ea5 : STD_LOGIC; 
  signal sig00000ea6 : STD_LOGIC; 
  signal sig00000ea7 : STD_LOGIC; 
  signal sig00000ea8 : STD_LOGIC; 
  signal sig00000ea9 : STD_LOGIC; 
  signal sig00000eaa : STD_LOGIC; 
  signal sig00000eab : STD_LOGIC; 
  signal sig00000eac : STD_LOGIC; 
  signal sig00000ead : STD_LOGIC; 
  signal sig00000eae : STD_LOGIC; 
  signal sig00000eaf : STD_LOGIC; 
  signal sig00000eb0 : STD_LOGIC; 
  signal sig00000eb1 : STD_LOGIC; 
  signal sig00000eb2 : STD_LOGIC; 
  signal sig00000eb3 : STD_LOGIC; 
  signal sig00000eb4 : STD_LOGIC; 
  signal sig00000eb5 : STD_LOGIC; 
  signal sig00000eb6 : STD_LOGIC; 
  signal sig00000eb7 : STD_LOGIC; 
  signal sig00000eb8 : STD_LOGIC; 
  signal sig00000eb9 : STD_LOGIC; 
  signal sig00000eba : STD_LOGIC; 
  signal sig00000ebb : STD_LOGIC; 
  signal sig00000ebc : STD_LOGIC; 
  signal sig00000ebd : STD_LOGIC; 
  signal sig00000ebe : STD_LOGIC; 
  signal sig00000ebf : STD_LOGIC; 
  signal sig00000ec0 : STD_LOGIC; 
  signal sig00000ec1 : STD_LOGIC; 
  signal sig00000ec2 : STD_LOGIC; 
  signal sig00000ec3 : STD_LOGIC; 
  signal sig00000ec4 : STD_LOGIC; 
  signal sig00000ec5 : STD_LOGIC; 
  signal sig00000ec6 : STD_LOGIC; 
  signal sig00000ec7 : STD_LOGIC; 
  signal sig00000ec8 : STD_LOGIC; 
  signal sig00000ec9 : STD_LOGIC; 
  signal sig00000eca : STD_LOGIC; 
  signal sig00000ecb : STD_LOGIC; 
  signal sig00000ecc : STD_LOGIC; 
  signal sig00000ecd : STD_LOGIC; 
  signal sig00000ece : STD_LOGIC; 
  signal sig00000ecf : STD_LOGIC; 
  signal sig00000ed0 : STD_LOGIC; 
  signal sig00000ed1 : STD_LOGIC; 
  signal sig00000ed2 : STD_LOGIC; 
  signal sig00000ed3 : STD_LOGIC; 
  signal sig00000ed4 : STD_LOGIC; 
  signal sig00000ed5 : STD_LOGIC; 
  signal sig00000ed6 : STD_LOGIC; 
  signal sig00000ed7 : STD_LOGIC; 
  signal sig00000ed8 : STD_LOGIC; 
  signal sig00000ed9 : STD_LOGIC; 
  signal sig00000eda : STD_LOGIC; 
  signal sig00000edb : STD_LOGIC; 
  signal sig00000edc : STD_LOGIC; 
  signal sig00000edd : STD_LOGIC; 
  signal sig00000ede : STD_LOGIC; 
  signal sig00000edf : STD_LOGIC; 
  signal sig00000ee0 : STD_LOGIC; 
  signal sig00000ee1 : STD_LOGIC; 
  signal sig00000ee2 : STD_LOGIC; 
  signal sig00000ee3 : STD_LOGIC; 
  signal sig00000ee4 : STD_LOGIC; 
  signal sig00000ee5 : STD_LOGIC; 
  signal sig00000ee6 : STD_LOGIC; 
  signal sig00000ee7 : STD_LOGIC; 
  signal sig00000ee8 : STD_LOGIC; 
  signal sig00000ee9 : STD_LOGIC; 
  signal sig00000eea : STD_LOGIC; 
  signal sig00000eeb : STD_LOGIC; 
  signal sig00000eec : STD_LOGIC; 
  signal sig00000eed : STD_LOGIC; 
  signal sig00000eee : STD_LOGIC; 
  signal sig00000eef : STD_LOGIC; 
  signal sig00000ef0 : STD_LOGIC; 
  signal sig00000ef1 : STD_LOGIC; 
  signal sig00000ef2 : STD_LOGIC; 
  signal sig00000ef3 : STD_LOGIC; 
  signal sig00000ef4 : STD_LOGIC; 
  signal sig00000ef5 : STD_LOGIC; 
  signal sig00000ef6 : STD_LOGIC; 
  signal sig00000ef7 : STD_LOGIC; 
  signal sig00000ef8 : STD_LOGIC; 
  signal sig00000ef9 : STD_LOGIC; 
  signal sig00000efa : STD_LOGIC; 
  signal sig00000efb : STD_LOGIC; 
  signal sig00000efc : STD_LOGIC; 
  signal sig00000efd : STD_LOGIC; 
  signal sig00000efe : STD_LOGIC; 
  signal sig00000eff : STD_LOGIC; 
  signal sig00000f00 : STD_LOGIC; 
  signal sig00000f01 : STD_LOGIC; 
  signal sig00000f02 : STD_LOGIC; 
  signal sig00000f03 : STD_LOGIC; 
  signal sig00000f04 : STD_LOGIC; 
  signal sig00000f05 : STD_LOGIC; 
  signal sig00000f06 : STD_LOGIC; 
  signal sig00000f07 : STD_LOGIC; 
  signal sig00000f08 : STD_LOGIC; 
  signal sig00000f09 : STD_LOGIC; 
  signal sig00000f0a : STD_LOGIC; 
  signal sig00000f0b : STD_LOGIC; 
  signal sig00000f0c : STD_LOGIC; 
  signal sig00000f0d : STD_LOGIC; 
  signal sig00000f0e : STD_LOGIC; 
  signal sig00000f0f : STD_LOGIC; 
  signal sig00000f10 : STD_LOGIC; 
  signal sig00000f11 : STD_LOGIC; 
  signal sig00000f12 : STD_LOGIC; 
  signal sig00000f13 : STD_LOGIC; 
  signal sig00000f14 : STD_LOGIC; 
  signal sig00000f15 : STD_LOGIC; 
  signal sig00000f16 : STD_LOGIC; 
  signal sig00000f17 : STD_LOGIC; 
  signal sig00000f18 : STD_LOGIC; 
  signal sig00000f19 : STD_LOGIC; 
  signal sig00000f1a : STD_LOGIC; 
  signal sig00000f1b : STD_LOGIC; 
  signal sig00000f1c : STD_LOGIC; 
  signal sig00000f1d : STD_LOGIC; 
  signal sig00000f1e : STD_LOGIC; 
  signal sig00000f1f : STD_LOGIC; 
  signal sig00000f20 : STD_LOGIC; 
  signal sig00000f21 : STD_LOGIC; 
  signal sig00000f22 : STD_LOGIC; 
  signal sig00000f23 : STD_LOGIC; 
  signal sig00000f24 : STD_LOGIC; 
  signal sig00000f25 : STD_LOGIC; 
  signal sig00000f26 : STD_LOGIC; 
  signal sig00000f27 : STD_LOGIC; 
  signal sig00000f28 : STD_LOGIC; 
  signal sig00000f29 : STD_LOGIC; 
  signal sig00000f2a : STD_LOGIC; 
  signal sig00000f2b : STD_LOGIC; 
  signal sig00000f2c : STD_LOGIC; 
  signal sig00000f2d : STD_LOGIC; 
  signal sig00000f2e : STD_LOGIC; 
  signal sig00000f2f : STD_LOGIC; 
  signal sig00000f30 : STD_LOGIC; 
  signal sig00000f31 : STD_LOGIC; 
  signal sig00000f32 : STD_LOGIC; 
  signal sig00000f33 : STD_LOGIC; 
  signal sig00000f34 : STD_LOGIC; 
  signal sig00000f35 : STD_LOGIC; 
  signal sig00000f36 : STD_LOGIC; 
  signal sig00000f37 : STD_LOGIC; 
  signal sig00000f38 : STD_LOGIC; 
  signal sig00000f39 : STD_LOGIC; 
  signal sig00000f3a : STD_LOGIC; 
  signal sig00000f3b : STD_LOGIC; 
  signal sig00000f3c : STD_LOGIC; 
  signal sig00000f3d : STD_LOGIC; 
  signal sig00000f3e : STD_LOGIC; 
  signal sig00000f3f : STD_LOGIC; 
  signal sig00000f40 : STD_LOGIC; 
  signal sig00000f41 : STD_LOGIC; 
  signal sig00000f42 : STD_LOGIC; 
  signal sig00000f43 : STD_LOGIC; 
  signal sig00000f44 : STD_LOGIC; 
  signal sig00000f45 : STD_LOGIC; 
  signal sig00000f46 : STD_LOGIC; 
  signal sig00000f47 : STD_LOGIC; 
  signal sig00000f48 : STD_LOGIC; 
  signal sig00000f49 : STD_LOGIC; 
  signal sig00000f4a : STD_LOGIC; 
  signal sig00000f4b : STD_LOGIC; 
  signal sig00000f4c : STD_LOGIC; 
  signal sig00000f4d : STD_LOGIC; 
  signal sig00000f4e : STD_LOGIC; 
  signal sig00000f4f : STD_LOGIC; 
  signal sig00000f50 : STD_LOGIC; 
  signal sig00000f51 : STD_LOGIC; 
  signal sig00000f52 : STD_LOGIC; 
  signal sig00000f53 : STD_LOGIC; 
  signal sig00000f54 : STD_LOGIC; 
  signal sig00000f55 : STD_LOGIC; 
  signal sig00000f56 : STD_LOGIC; 
  signal sig00000f57 : STD_LOGIC; 
  signal sig00000f58 : STD_LOGIC; 
  signal sig00000f59 : STD_LOGIC; 
  signal sig00000f5a : STD_LOGIC; 
  signal sig00000f5b : STD_LOGIC; 
  signal sig00000f5c : STD_LOGIC; 
  signal sig00000f5d : STD_LOGIC; 
  signal sig00000f5e : STD_LOGIC; 
  signal sig00000f5f : STD_LOGIC; 
  signal sig00000f60 : STD_LOGIC; 
  signal sig00000f61 : STD_LOGIC; 
  signal sig00000f62 : STD_LOGIC; 
  signal sig00000f63 : STD_LOGIC; 
  signal sig00000f64 : STD_LOGIC; 
  signal sig00000f65 : STD_LOGIC; 
  signal sig00000f66 : STD_LOGIC; 
  signal sig00000f67 : STD_LOGIC; 
  signal sig00000f68 : STD_LOGIC; 
  signal sig00000f69 : STD_LOGIC; 
  signal sig00000f6a : STD_LOGIC; 
  signal sig00000f6b : STD_LOGIC; 
  signal sig00000f6c : STD_LOGIC; 
  signal sig00000f6d : STD_LOGIC; 
  signal sig00000f6e : STD_LOGIC; 
  signal sig00000f6f : STD_LOGIC; 
  signal sig00000f70 : STD_LOGIC; 
  signal sig00000f71 : STD_LOGIC; 
  signal sig00000f72 : STD_LOGIC; 
  signal sig00000f73 : STD_LOGIC; 
  signal sig00000f74 : STD_LOGIC; 
  signal sig00000f75 : STD_LOGIC; 
  signal sig00000f76 : STD_LOGIC; 
  signal sig00000f77 : STD_LOGIC; 
  signal sig00000f78 : STD_LOGIC; 
  signal sig00000f79 : STD_LOGIC; 
  signal sig00000f7a : STD_LOGIC; 
  signal sig00000f7b : STD_LOGIC; 
  signal sig00000f7c : STD_LOGIC; 
  signal sig00000f7d : STD_LOGIC; 
  signal sig00000f7e : STD_LOGIC; 
  signal sig00000f7f : STD_LOGIC; 
  signal sig00000f80 : STD_LOGIC; 
  signal sig00000f81 : STD_LOGIC; 
  signal sig00000f82 : STD_LOGIC; 
  signal sig00000f83 : STD_LOGIC; 
  signal sig00000f84 : STD_LOGIC; 
  signal sig00000f85 : STD_LOGIC; 
  signal sig00000f86 : STD_LOGIC; 
  signal sig00000f87 : STD_LOGIC; 
  signal sig00000f88 : STD_LOGIC; 
  signal sig00000f89 : STD_LOGIC; 
  signal sig00000f8a : STD_LOGIC; 
  signal sig00000f8b : STD_LOGIC; 
  signal sig00000f8c : STD_LOGIC; 
  signal sig00000f8d : STD_LOGIC; 
  signal sig00000f8e : STD_LOGIC; 
  signal sig00000f8f : STD_LOGIC; 
  signal sig00000f90 : STD_LOGIC; 
  signal sig00000f91 : STD_LOGIC; 
  signal sig00000f92 : STD_LOGIC; 
  signal sig00000f93 : STD_LOGIC; 
  signal sig00000f94 : STD_LOGIC; 
  signal sig00000f95 : STD_LOGIC; 
  signal sig00000f96 : STD_LOGIC; 
  signal sig00000f97 : STD_LOGIC; 
  signal sig00000f98 : STD_LOGIC; 
  signal blk00000065_blk00000066_sig00000fdb : STD_LOGIC; 
  signal blk00000065_blk00000066_sig00000fda : STD_LOGIC; 
  signal blk00000065_blk00000066_sig00000fd9 : STD_LOGIC; 
  signal blk00000065_blk00000066_sig00000fd8 : STD_LOGIC; 
  signal blk00000065_blk00000066_sig00000fd7 : STD_LOGIC; 
  signal blk00000065_blk00000066_sig00000fd6 : STD_LOGIC; 
  signal blk00000065_blk00000066_sig00000fd5 : STD_LOGIC; 
  signal blk00000065_blk00000066_sig00000fd4 : STD_LOGIC; 
  signal blk00000065_blk00000066_sig00000fd3 : STD_LOGIC; 
  signal blk00000065_blk00000066_sig00000fd2 : STD_LOGIC; 
  signal blk00000065_blk00000066_sig00000fd1 : STD_LOGIC; 
  signal blk00000065_blk00000066_sig00000fd0 : STD_LOGIC; 
  signal blk00000065_blk00000066_sig00000fcf : STD_LOGIC; 
  signal blk00000065_blk00000066_sig00000fce : STD_LOGIC; 
  signal blk00000081_blk00000082_sig0000101e : STD_LOGIC; 
  signal blk00000081_blk00000082_sig0000101d : STD_LOGIC; 
  signal blk00000081_blk00000082_sig0000101c : STD_LOGIC; 
  signal blk00000081_blk00000082_sig0000101b : STD_LOGIC; 
  signal blk00000081_blk00000082_sig0000101a : STD_LOGIC; 
  signal blk00000081_blk00000082_sig00001019 : STD_LOGIC; 
  signal blk00000081_blk00000082_sig00001018 : STD_LOGIC; 
  signal blk00000081_blk00000082_sig00001017 : STD_LOGIC; 
  signal blk00000081_blk00000082_sig00001016 : STD_LOGIC; 
  signal blk00000081_blk00000082_sig00001015 : STD_LOGIC; 
  signal blk00000081_blk00000082_sig00001014 : STD_LOGIC; 
  signal blk00000081_blk00000082_sig00001013 : STD_LOGIC; 
  signal blk00000081_blk00000082_sig00001012 : STD_LOGIC; 
  signal blk00000081_blk00000082_sig00001011 : STD_LOGIC; 
  signal blk000000ed_sig0000103e : STD_LOGIC; 
  signal blk000000ed_sig0000103d : STD_LOGIC; 
  signal blk000000ed_sig0000103c : STD_LOGIC; 
  signal blk000000ed_sig0000103b : STD_LOGIC; 
  signal blk000000ed_sig0000103a : STD_LOGIC; 
  signal blk000000ed_sig00001039 : STD_LOGIC; 
  signal blk000000ed_sig00001038 : STD_LOGIC; 
  signal blk000000ed_sig00001037 : STD_LOGIC; 
  signal blk000000ed_sig00001036 : STD_LOGIC; 
  signal blk000000ed_sig00001035 : STD_LOGIC; 
  signal blk000000ed_sig00001034 : STD_LOGIC; 
  signal blk000000ed_sig00001033 : STD_LOGIC; 
  signal blk000000ed_sig00001032 : STD_LOGIC; 
  signal blk000000ed_sig00001031 : STD_LOGIC; 
  signal blk000000ed_sig00001030 : STD_LOGIC; 
  signal blk000000ed_sig0000102f : STD_LOGIC; 
  signal blk00000104_sig0000105e : STD_LOGIC; 
  signal blk00000104_sig0000105d : STD_LOGIC; 
  signal blk00000104_sig0000105c : STD_LOGIC; 
  signal blk00000104_sig0000105b : STD_LOGIC; 
  signal blk00000104_sig0000105a : STD_LOGIC; 
  signal blk00000104_sig00001059 : STD_LOGIC; 
  signal blk00000104_sig00001058 : STD_LOGIC; 
  signal blk00000104_sig00001057 : STD_LOGIC; 
  signal blk00000104_sig00001056 : STD_LOGIC; 
  signal blk00000104_sig00001055 : STD_LOGIC; 
  signal blk00000104_sig00001054 : STD_LOGIC; 
  signal blk00000104_sig00001053 : STD_LOGIC; 
  signal blk00000104_sig00001052 : STD_LOGIC; 
  signal blk00000104_sig00001051 : STD_LOGIC; 
  signal blk00000104_sig00001050 : STD_LOGIC; 
  signal blk00000104_sig0000104f : STD_LOGIC; 
  signal blk0000011b_sig0000107e : STD_LOGIC; 
  signal blk0000011b_sig0000107d : STD_LOGIC; 
  signal blk0000011b_sig0000107c : STD_LOGIC; 
  signal blk0000011b_sig0000107b : STD_LOGIC; 
  signal blk0000011b_sig0000107a : STD_LOGIC; 
  signal blk0000011b_sig00001079 : STD_LOGIC; 
  signal blk0000011b_sig00001078 : STD_LOGIC; 
  signal blk0000011b_sig00001077 : STD_LOGIC; 
  signal blk0000011b_sig00001076 : STD_LOGIC; 
  signal blk0000011b_sig00001075 : STD_LOGIC; 
  signal blk0000011b_sig00001074 : STD_LOGIC; 
  signal blk0000011b_sig00001073 : STD_LOGIC; 
  signal blk0000011b_sig00001072 : STD_LOGIC; 
  signal blk0000011b_sig00001071 : STD_LOGIC; 
  signal blk0000011b_sig00001070 : STD_LOGIC; 
  signal blk0000011b_sig0000106f : STD_LOGIC; 
  signal blk0000014b_sig0000109e : STD_LOGIC; 
  signal blk0000014b_sig0000109d : STD_LOGIC; 
  signal blk0000014b_sig0000109c : STD_LOGIC; 
  signal blk0000014b_sig0000109b : STD_LOGIC; 
  signal blk0000014b_sig0000109a : STD_LOGIC; 
  signal blk0000014b_sig00001099 : STD_LOGIC; 
  signal blk0000014b_sig00001098 : STD_LOGIC; 
  signal blk0000014b_sig00001097 : STD_LOGIC; 
  signal blk0000014b_sig00001096 : STD_LOGIC; 
  signal blk0000014b_sig00001095 : STD_LOGIC; 
  signal blk0000014b_sig00001094 : STD_LOGIC; 
  signal blk0000014b_sig00001093 : STD_LOGIC; 
  signal blk0000014b_sig00001092 : STD_LOGIC; 
  signal blk0000014b_sig00001091 : STD_LOGIC; 
  signal blk0000014b_sig00001090 : STD_LOGIC; 
  signal blk0000014b_sig0000108f : STD_LOGIC; 
  signal blk0000017b_blk0000017c_sig000010b0 : STD_LOGIC; 
  signal blk0000017b_blk0000017c_sig000010af : STD_LOGIC; 
  signal blk0000017b_blk0000017c_sig000010ae : STD_LOGIC; 
  signal blk00000181_blk00000182_sig000010c2 : STD_LOGIC; 
  signal blk00000181_blk00000182_sig000010c1 : STD_LOGIC; 
  signal blk00000181_blk00000182_sig000010c0 : STD_LOGIC; 
  signal blk00000187_blk00000188_sig000010d4 : STD_LOGIC; 
  signal blk00000187_blk00000188_sig000010d3 : STD_LOGIC; 
  signal blk00000187_blk00000188_sig000010d2 : STD_LOGIC; 
  signal blk0000018d_sig000010e3 : STD_LOGIC; 
  signal blk0000018d_sig000010e2 : STD_LOGIC; 
  signal blk0000018d_sig000010e1 : STD_LOGIC; 
  signal blk0000018d_sig000010e0 : STD_LOGIC; 
  signal blk0000018d_sig000010df : STD_LOGIC; 
  signal blk0000018d_blk0000018e_sig000010ea : STD_LOGIC; 
  signal blk0000018d_blk0000018e_sig000010e9 : STD_LOGIC; 
  signal blk0000018d_blk0000018e_sig000010e8 : STD_LOGIC; 
  signal blk00000193_sig000010f9 : STD_LOGIC; 
  signal blk00000193_sig000010f8 : STD_LOGIC; 
  signal blk00000193_sig000010f7 : STD_LOGIC; 
  signal blk00000193_sig000010f6 : STD_LOGIC; 
  signal blk00000193_blk00000194_sig00001103 : STD_LOGIC; 
  signal blk00000193_blk00000194_sig00001102 : STD_LOGIC; 
  signal blk00000193_blk00000194_sig00001101 : STD_LOGIC; 
  signal blk00000193_blk00000194_sig00001100 : STD_LOGIC; 
  signal blk000001aa_sig00001123 : STD_LOGIC; 
  signal blk000001aa_sig00001122 : STD_LOGIC; 
  signal blk000001aa_sig00001121 : STD_LOGIC; 
  signal blk000001aa_sig00001120 : STD_LOGIC; 
  signal blk000001aa_sig0000111f : STD_LOGIC; 
  signal blk000001aa_sig0000111e : STD_LOGIC; 
  signal blk000001aa_sig0000111d : STD_LOGIC; 
  signal blk000001aa_sig0000111c : STD_LOGIC; 
  signal blk000001aa_sig0000111b : STD_LOGIC; 
  signal blk000001aa_sig0000111a : STD_LOGIC; 
  signal blk000001aa_sig00001119 : STD_LOGIC; 
  signal blk000001aa_sig00001118 : STD_LOGIC; 
  signal blk000001aa_sig00001117 : STD_LOGIC; 
  signal blk000001aa_sig00001116 : STD_LOGIC; 
  signal blk000001aa_sig00001115 : STD_LOGIC; 
  signal blk000001aa_sig00001114 : STD_LOGIC; 
  signal blk000001d2_sig00001143 : STD_LOGIC; 
  signal blk000001d2_sig00001142 : STD_LOGIC; 
  signal blk000001d2_sig00001141 : STD_LOGIC; 
  signal blk000001d2_sig00001140 : STD_LOGIC; 
  signal blk000001d2_sig0000113f : STD_LOGIC; 
  signal blk000001d2_sig0000113e : STD_LOGIC; 
  signal blk000001d2_sig0000113d : STD_LOGIC; 
  signal blk000001d2_sig0000113c : STD_LOGIC; 
  signal blk000001d2_sig0000113b : STD_LOGIC; 
  signal blk000001d2_sig0000113a : STD_LOGIC; 
  signal blk000001d2_sig00001139 : STD_LOGIC; 
  signal blk000001d2_sig00001138 : STD_LOGIC; 
  signal blk000001d2_sig00001137 : STD_LOGIC; 
  signal blk000001d2_sig00001136 : STD_LOGIC; 
  signal blk000001d2_sig00001135 : STD_LOGIC; 
  signal blk000001d2_sig00001134 : STD_LOGIC; 
  signal blk000001fa_blk000001fb_sig00001155 : STD_LOGIC; 
  signal blk000001fa_blk000001fb_sig00001154 : STD_LOGIC; 
  signal blk000001fa_blk000001fb_sig00001153 : STD_LOGIC; 
  signal blk00000200_blk00000201_sig00001198 : STD_LOGIC; 
  signal blk00000200_blk00000201_sig00001197 : STD_LOGIC; 
  signal blk00000200_blk00000201_sig00001196 : STD_LOGIC; 
  signal blk00000200_blk00000201_sig00001195 : STD_LOGIC; 
  signal blk00000200_blk00000201_sig00001194 : STD_LOGIC; 
  signal blk00000200_blk00000201_sig00001193 : STD_LOGIC; 
  signal blk00000200_blk00000201_sig00001192 : STD_LOGIC; 
  signal blk00000200_blk00000201_sig00001191 : STD_LOGIC; 
  signal blk00000200_blk00000201_sig00001190 : STD_LOGIC; 
  signal blk00000200_blk00000201_sig0000118f : STD_LOGIC; 
  signal blk00000200_blk00000201_sig0000118e : STD_LOGIC; 
  signal blk00000200_blk00000201_sig0000118d : STD_LOGIC; 
  signal blk00000200_blk00000201_sig0000118c : STD_LOGIC; 
  signal blk00000200_blk00000201_sig0000118b : STD_LOGIC; 
  signal blk0000021c_blk0000021d_sig000011db : STD_LOGIC; 
  signal blk0000021c_blk0000021d_sig000011da : STD_LOGIC; 
  signal blk0000021c_blk0000021d_sig000011d9 : STD_LOGIC; 
  signal blk0000021c_blk0000021d_sig000011d8 : STD_LOGIC; 
  signal blk0000021c_blk0000021d_sig000011d7 : STD_LOGIC; 
  signal blk0000021c_blk0000021d_sig000011d6 : STD_LOGIC; 
  signal blk0000021c_blk0000021d_sig000011d5 : STD_LOGIC; 
  signal blk0000021c_blk0000021d_sig000011d4 : STD_LOGIC; 
  signal blk0000021c_blk0000021d_sig000011d3 : STD_LOGIC; 
  signal blk0000021c_blk0000021d_sig000011d2 : STD_LOGIC; 
  signal blk0000021c_blk0000021d_sig000011d1 : STD_LOGIC; 
  signal blk0000021c_blk0000021d_sig000011d0 : STD_LOGIC; 
  signal blk0000021c_blk0000021d_sig000011cf : STD_LOGIC; 
  signal blk0000021c_blk0000021d_sig000011ce : STD_LOGIC; 
  signal blk00000287_blk00000288_sig00001263 : STD_LOGIC; 
  signal blk00000287_blk00000288_sig00001262 : STD_LOGIC; 
  signal blk00000287_blk00000288_sig00001261 : STD_LOGIC; 
  signal blk00000287_blk00000288_sig00001260 : STD_LOGIC; 
  signal blk00000287_blk00000288_sig0000125f : STD_LOGIC; 
  signal blk00000287_blk00000288_sig0000125e : STD_LOGIC; 
  signal blk00000287_blk00000288_sig0000125d : STD_LOGIC; 
  signal blk00000287_blk00000288_sig0000125c : STD_LOGIC; 
  signal blk00000287_blk00000288_sig0000125b : STD_LOGIC; 
  signal blk00000287_blk00000288_sig0000125a : STD_LOGIC; 
  signal blk00000287_blk00000288_sig00001259 : STD_LOGIC; 
  signal blk00000287_blk00000288_sig00001258 : STD_LOGIC; 
  signal blk00000287_blk00000288_sig00001257 : STD_LOGIC; 
  signal blk00000287_blk00000288_sig00001256 : STD_LOGIC; 
  signal blk00000287_blk00000288_sig00001255 : STD_LOGIC; 
  signal blk00000287_blk00000288_sig00001254 : STD_LOGIC; 
  signal blk00000287_blk00000288_sig00001253 : STD_LOGIC; 
  signal blk00000287_blk00000288_sig00001252 : STD_LOGIC; 
  signal blk00000287_blk00000288_sig00001251 : STD_LOGIC; 
  signal blk00000287_blk00000288_sig00001250 : STD_LOGIC; 
  signal blk00000287_blk00000288_sig0000124f : STD_LOGIC; 
  signal blk00000287_blk00000288_sig0000124e : STD_LOGIC; 
  signal blk00000287_blk00000288_sig0000124d : STD_LOGIC; 
  signal blk00000287_blk00000288_sig0000124c : STD_LOGIC; 
  signal blk00000287_blk00000288_sig0000124b : STD_LOGIC; 
  signal blk00000287_blk00000288_sig0000124a : STD_LOGIC; 
  signal blk00000287_blk00000288_sig00001249 : STD_LOGIC; 
  signal blk00000287_blk00000288_sig00001248 : STD_LOGIC; 
  signal blk000002bf_sig000012b8 : STD_LOGIC; 
  signal blk000002bf_sig000012b7 : STD_LOGIC; 
  signal blk000002bf_sig000012b6 : STD_LOGIC; 
  signal blk000002bf_sig000012b5 : STD_LOGIC; 
  signal blk000002bf_sig000012b4 : STD_LOGIC; 
  signal blk000002bf_sig000012b3 : STD_LOGIC; 
  signal blk000002bf_sig000012b2 : STD_LOGIC; 
  signal blk000002bf_sig000012b1 : STD_LOGIC; 
  signal blk000002bf_sig000012b0 : STD_LOGIC; 
  signal blk000002bf_sig000012af : STD_LOGIC; 
  signal blk000002bf_sig000012ae : STD_LOGIC; 
  signal blk000002bf_sig000012ad : STD_LOGIC; 
  signal blk000002bf_sig000012ac : STD_LOGIC; 
  signal blk000002bf_sig000012ab : STD_LOGIC; 
  signal blk000002bf_sig000012aa : STD_LOGIC; 
  signal blk000002bf_sig000012a9 : STD_LOGIC; 
  signal blk000002bf_sig000012a8 : STD_LOGIC; 
  signal blk000002bf_sig000012a7 : STD_LOGIC; 
  signal blk000002bf_sig000012a6 : STD_LOGIC; 
  signal blk000002bf_sig000012a5 : STD_LOGIC; 
  signal blk000002bf_sig000012a4 : STD_LOGIC; 
  signal blk000002bf_sig000012a3 : STD_LOGIC; 
  signal blk000002bf_sig000012a2 : STD_LOGIC; 
  signal blk000002bf_sig000012a1 : STD_LOGIC; 
  signal blk000002bf_sig000012a0 : STD_LOGIC; 
  signal blk000002bf_sig0000129f : STD_LOGIC; 
  signal blk000002bf_sig0000129e : STD_LOGIC; 
  signal blk000002bf_sig0000129d : STD_LOGIC; 
  signal blk000002bf_sig0000129c : STD_LOGIC; 
  signal blk000002bf_sig0000129b : STD_LOGIC; 
  signal blk000002bf_sig0000129a : STD_LOGIC; 
  signal blk000002bf_sig00001299 : STD_LOGIC; 
  signal blk000002bf_sig00001298 : STD_LOGIC; 
  signal blk000002bf_sig00001297 : STD_LOGIC; 
  signal blk000002bf_sig00001296 : STD_LOGIC; 
  signal blk000002bf_sig00001295 : STD_LOGIC; 
  signal blk000002bf_sig00001294 : STD_LOGIC; 
  signal blk000002bf_sig00001293 : STD_LOGIC; 
  signal blk000002bf_sig00001292 : STD_LOGIC; 
  signal blk000002bf_sig00001291 : STD_LOGIC; 
  signal blk000002bf_sig00001290 : STD_LOGIC; 
  signal blk000002bf_sig0000128f : STD_LOGIC; 
  signal blk000002f8_sig0000130d : STD_LOGIC; 
  signal blk000002f8_sig0000130c : STD_LOGIC; 
  signal blk000002f8_sig0000130b : STD_LOGIC; 
  signal blk000002f8_sig0000130a : STD_LOGIC; 
  signal blk000002f8_sig00001309 : STD_LOGIC; 
  signal blk000002f8_sig00001308 : STD_LOGIC; 
  signal blk000002f8_sig00001307 : STD_LOGIC; 
  signal blk000002f8_sig00001306 : STD_LOGIC; 
  signal blk000002f8_sig00001305 : STD_LOGIC; 
  signal blk000002f8_sig00001304 : STD_LOGIC; 
  signal blk000002f8_sig00001303 : STD_LOGIC; 
  signal blk000002f8_sig00001302 : STD_LOGIC; 
  signal blk000002f8_sig00001301 : STD_LOGIC; 
  signal blk000002f8_sig00001300 : STD_LOGIC; 
  signal blk000002f8_sig000012ff : STD_LOGIC; 
  signal blk000002f8_sig000012fe : STD_LOGIC; 
  signal blk000002f8_sig000012fd : STD_LOGIC; 
  signal blk000002f8_sig000012fc : STD_LOGIC; 
  signal blk000002f8_sig000012fb : STD_LOGIC; 
  signal blk000002f8_sig000012fa : STD_LOGIC; 
  signal blk000002f8_sig000012f9 : STD_LOGIC; 
  signal blk000002f8_sig000012f8 : STD_LOGIC; 
  signal blk000002f8_sig000012f7 : STD_LOGIC; 
  signal blk000002f8_sig000012f6 : STD_LOGIC; 
  signal blk000002f8_sig000012f5 : STD_LOGIC; 
  signal blk000002f8_sig000012f4 : STD_LOGIC; 
  signal blk000002f8_sig000012f3 : STD_LOGIC; 
  signal blk000002f8_sig000012f2 : STD_LOGIC; 
  signal blk000002f8_sig000012f1 : STD_LOGIC; 
  signal blk000002f8_sig000012f0 : STD_LOGIC; 
  signal blk000002f8_sig000012ef : STD_LOGIC; 
  signal blk000002f8_sig000012ee : STD_LOGIC; 
  signal blk000002f8_sig000012ed : STD_LOGIC; 
  signal blk000002f8_sig000012ec : STD_LOGIC; 
  signal blk000002f8_sig000012eb : STD_LOGIC; 
  signal blk000002f8_sig000012ea : STD_LOGIC; 
  signal blk000002f8_sig000012e9 : STD_LOGIC; 
  signal blk000002f8_sig000012e8 : STD_LOGIC; 
  signal blk000002f8_sig000012e7 : STD_LOGIC; 
  signal blk000002f8_sig000012e6 : STD_LOGIC; 
  signal blk000002f8_sig000012e5 : STD_LOGIC; 
  signal blk000002f8_sig000012e4 : STD_LOGIC; 
  signal blk00000331_sig0000136e : STD_LOGIC; 
  signal blk00000331_sig0000136d : STD_LOGIC; 
  signal blk00000331_sig0000136c : STD_LOGIC; 
  signal blk00000331_sig0000136b : STD_LOGIC; 
  signal blk00000331_sig0000136a : STD_LOGIC; 
  signal blk00000331_sig00001369 : STD_LOGIC; 
  signal blk00000331_sig00001368 : STD_LOGIC; 
  signal blk00000331_sig00001367 : STD_LOGIC; 
  signal blk00000331_sig00001366 : STD_LOGIC; 
  signal blk00000331_sig00001365 : STD_LOGIC; 
  signal blk00000331_sig00001364 : STD_LOGIC; 
  signal blk00000331_sig00001363 : STD_LOGIC; 
  signal blk00000331_sig00001362 : STD_LOGIC; 
  signal blk00000331_sig00001361 : STD_LOGIC; 
  signal blk00000331_sig00001360 : STD_LOGIC; 
  signal blk00000331_sig0000135f : STD_LOGIC; 
  signal blk00000331_sig0000135e : STD_LOGIC; 
  signal blk00000331_sig0000135d : STD_LOGIC; 
  signal blk00000331_sig0000135c : STD_LOGIC; 
  signal blk00000331_sig0000135b : STD_LOGIC; 
  signal blk00000331_sig0000135a : STD_LOGIC; 
  signal blk00000331_sig00001359 : STD_LOGIC; 
  signal blk00000331_sig00001358 : STD_LOGIC; 
  signal blk00000331_sig00001357 : STD_LOGIC; 
  signal blk00000331_sig00001356 : STD_LOGIC; 
  signal blk00000331_sig00001355 : STD_LOGIC; 
  signal blk00000331_sig00001354 : STD_LOGIC; 
  signal blk00000331_sig00001353 : STD_LOGIC; 
  signal blk00000331_sig00001352 : STD_LOGIC; 
  signal blk00000331_sig00001351 : STD_LOGIC; 
  signal blk00000331_sig00001350 : STD_LOGIC; 
  signal blk00000331_sig0000134f : STD_LOGIC; 
  signal blk00000331_sig0000134e : STD_LOGIC; 
  signal blk00000331_sig0000134d : STD_LOGIC; 
  signal blk00000331_sig0000134c : STD_LOGIC; 
  signal blk00000331_sig0000134b : STD_LOGIC; 
  signal blk00000331_sig0000134a : STD_LOGIC; 
  signal blk00000331_sig00001349 : STD_LOGIC; 
  signal blk00000331_sig00001348 : STD_LOGIC; 
  signal blk00000331_sig00001347 : STD_LOGIC; 
  signal blk00000331_sig00001346 : STD_LOGIC; 
  signal blk00000331_sig00001345 : STD_LOGIC; 
  signal blk00000331_sig00001344 : STD_LOGIC; 
  signal blk00000331_sig00001343 : STD_LOGIC; 
  signal blk00000331_sig00001342 : STD_LOGIC; 
  signal blk00000331_sig00001341 : STD_LOGIC; 
  signal blk00000331_sig00001340 : STD_LOGIC; 
  signal blk00000331_sig0000133f : STD_LOGIC; 
  signal blk00000331_sig0000133e : STD_LOGIC; 
  signal blk00000331_sig0000133d : STD_LOGIC; 
  signal blk00000331_sig0000133c : STD_LOGIC; 
  signal blk00000331_sig0000133b : STD_LOGIC; 
  signal blk00000331_sig0000133a : STD_LOGIC; 
  signal blk00000331_sig00001339 : STD_LOGIC; 
  signal blk00000376_sig000013cf : STD_LOGIC; 
  signal blk00000376_sig000013ce : STD_LOGIC; 
  signal blk00000376_sig000013cd : STD_LOGIC; 
  signal blk00000376_sig000013cc : STD_LOGIC; 
  signal blk00000376_sig000013cb : STD_LOGIC; 
  signal blk00000376_sig000013ca : STD_LOGIC; 
  signal blk00000376_sig000013c9 : STD_LOGIC; 
  signal blk00000376_sig000013c8 : STD_LOGIC; 
  signal blk00000376_sig000013c7 : STD_LOGIC; 
  signal blk00000376_sig000013c6 : STD_LOGIC; 
  signal blk00000376_sig000013c5 : STD_LOGIC; 
  signal blk00000376_sig000013c4 : STD_LOGIC; 
  signal blk00000376_sig000013c3 : STD_LOGIC; 
  signal blk00000376_sig000013c2 : STD_LOGIC; 
  signal blk00000376_sig000013c1 : STD_LOGIC; 
  signal blk00000376_sig000013c0 : STD_LOGIC; 
  signal blk00000376_sig000013bf : STD_LOGIC; 
  signal blk00000376_sig000013be : STD_LOGIC; 
  signal blk00000376_sig000013bd : STD_LOGIC; 
  signal blk00000376_sig000013bc : STD_LOGIC; 
  signal blk00000376_sig000013bb : STD_LOGIC; 
  signal blk00000376_sig000013ba : STD_LOGIC; 
  signal blk00000376_sig000013b9 : STD_LOGIC; 
  signal blk00000376_sig000013b8 : STD_LOGIC; 
  signal blk00000376_sig000013b7 : STD_LOGIC; 
  signal blk00000376_sig000013b6 : STD_LOGIC; 
  signal blk00000376_sig000013b5 : STD_LOGIC; 
  signal blk00000376_sig000013b4 : STD_LOGIC; 
  signal blk00000376_sig000013b3 : STD_LOGIC; 
  signal blk00000376_sig000013b2 : STD_LOGIC; 
  signal blk00000376_sig000013b1 : STD_LOGIC; 
  signal blk00000376_sig000013b0 : STD_LOGIC; 
  signal blk00000376_sig000013af : STD_LOGIC; 
  signal blk00000376_sig000013ae : STD_LOGIC; 
  signal blk00000376_sig000013ad : STD_LOGIC; 
  signal blk00000376_sig000013ac : STD_LOGIC; 
  signal blk00000376_sig000013ab : STD_LOGIC; 
  signal blk00000376_sig000013aa : STD_LOGIC; 
  signal blk00000376_sig000013a9 : STD_LOGIC; 
  signal blk00000376_sig000013a8 : STD_LOGIC; 
  signal blk00000376_sig000013a7 : STD_LOGIC; 
  signal blk00000376_sig000013a6 : STD_LOGIC; 
  signal blk00000376_sig000013a5 : STD_LOGIC; 
  signal blk00000376_sig000013a4 : STD_LOGIC; 
  signal blk00000376_sig000013a3 : STD_LOGIC; 
  signal blk00000376_sig000013a2 : STD_LOGIC; 
  signal blk00000376_sig000013a1 : STD_LOGIC; 
  signal blk00000376_sig000013a0 : STD_LOGIC; 
  signal blk00000376_sig0000139f : STD_LOGIC; 
  signal blk00000376_sig0000139e : STD_LOGIC; 
  signal blk00000376_sig0000139d : STD_LOGIC; 
  signal blk00000376_sig0000139c : STD_LOGIC; 
  signal blk00000376_sig0000139b : STD_LOGIC; 
  signal blk00000376_sig0000139a : STD_LOGIC; 
  signal blk000003bb_sig000013de : STD_LOGIC; 
  signal blk000003bb_sig000013dd : STD_LOGIC; 
  signal blk000003bb_sig000013dc : STD_LOGIC; 
  signal blk000003bb_sig000013da : STD_LOGIC; 
  signal blk000003bb_sig000013d9 : STD_LOGIC; 
  signal blk000003bb_blk000003bc_sig000013e4 : STD_LOGIC; 
  signal blk000003bb_blk000003bc_sig000013e3 : STD_LOGIC; 
  signal blk000003c0_blk000003c1_sig00001408 : STD_LOGIC; 
  signal blk000003c0_blk000003c1_sig00001407 : STD_LOGIC; 
  signal blk000003c0_blk000003c1_sig00001406 : STD_LOGIC; 
  signal blk000003c0_blk000003c1_sig00001405 : STD_LOGIC; 
  signal blk000003c0_blk000003c1_sig00001404 : STD_LOGIC; 
  signal blk000003c0_blk000003c1_sig00001403 : STD_LOGIC; 
  signal blk000003c0_blk000003c1_sig00001402 : STD_LOGIC; 
  signal blk000003cf_blk000003d0_sig00001413 : STD_LOGIC; 
  signal blk000003cf_blk000003d0_sig00001412 : STD_LOGIC; 
  signal blk000003cf_blk000003d0_sig00001411 : STD_LOGIC; 
  signal blk000003d5_blk000003d6_sig0000141f : STD_LOGIC; 
  signal blk000003d5_blk000003d6_sig0000141e : STD_LOGIC; 
  signal blk000003d5_blk000003d6_sig0000141d : STD_LOGIC; 
  signal blk000003db_blk000003dc_sig00001429 : STD_LOGIC; 
  signal blk000003db_blk000003dc_sig00001428 : STD_LOGIC; 
  signal blk000003e0_blk000003e1_sig00001439 : STD_LOGIC; 
  signal blk000003e0_blk000003e1_sig00001438 : STD_LOGIC; 
  signal blk000003e0_blk000003e1_sig00001437 : STD_LOGIC; 
  signal blk000003e0_blk000003e1_sig00001436 : STD_LOGIC; 
  signal blk000003e8_blk000003e9_sig00001452 : STD_LOGIC; 
  signal blk000003e8_blk000003e9_sig00001451 : STD_LOGIC; 
  signal blk000003e8_blk000003e9_sig00001450 : STD_LOGIC; 
  signal blk000003e8_blk000003e9_sig0000144f : STD_LOGIC; 
  signal blk000003e8_blk000003e9_sig0000144e : STD_LOGIC; 
  signal blk000004a0_blk000004a1_sig00001463 : STD_LOGIC; 
  signal blk000004a0_blk000004a1_sig00001462 : STD_LOGIC; 
  signal blk000004a5_blk000004a6_sig00001474 : STD_LOGIC; 
  signal blk000004a5_blk000004a6_sig00001473 : STD_LOGIC; 
  signal blk000004aa_blk000004ab_sig00001485 : STD_LOGIC; 
  signal blk000004aa_blk000004ab_sig00001484 : STD_LOGIC; 
  signal blk000004af_blk000004b0_sig00001496 : STD_LOGIC; 
  signal blk000004af_blk000004b0_sig00001495 : STD_LOGIC; 
  signal blk000004b4_blk000004b5_sig000014a2 : STD_LOGIC; 
  signal blk000004b4_blk000004b5_sig000014a1 : STD_LOGIC; 
  signal blk000004b4_blk000004b5_sig000014a0 : STD_LOGIC; 
  signal blk000004ba_blk000004bb_sig000014ef : STD_LOGIC; 
  signal blk000004ba_blk000004bb_sig000014ee : STD_LOGIC; 
  signal blk000004ba_blk000004bb_sig000014ed : STD_LOGIC; 
  signal blk000004ba_blk000004bb_sig000014ec : STD_LOGIC; 
  signal blk000004ba_blk000004bb_sig000014eb : STD_LOGIC; 
  signal blk000004ba_blk000004bb_sig000014ea : STD_LOGIC; 
  signal blk000004ba_blk000004bb_sig000014e9 : STD_LOGIC; 
  signal blk000004ba_blk000004bb_sig000014e8 : STD_LOGIC; 
  signal blk000004ba_blk000004bb_sig000014e7 : STD_LOGIC; 
  signal blk000004ba_blk000004bb_sig000014e6 : STD_LOGIC; 
  signal blk000004ba_blk000004bb_sig000014e5 : STD_LOGIC; 
  signal blk000004ba_blk000004bb_sig000014e4 : STD_LOGIC; 
  signal blk000004ba_blk000004bb_sig000014e3 : STD_LOGIC; 
  signal blk000004ba_blk000004bb_sig000014e2 : STD_LOGIC; 
  signal blk000004ba_blk000004bb_sig000014e1 : STD_LOGIC; 
  signal blk000004ba_blk000004bb_sig000014e0 : STD_LOGIC; 
  signal blk000004da_blk000004db_sig0000153c : STD_LOGIC; 
  signal blk000004da_blk000004db_sig0000153b : STD_LOGIC; 
  signal blk000004da_blk000004db_sig0000153a : STD_LOGIC; 
  signal blk000004da_blk000004db_sig00001539 : STD_LOGIC; 
  signal blk000004da_blk000004db_sig00001538 : STD_LOGIC; 
  signal blk000004da_blk000004db_sig00001537 : STD_LOGIC; 
  signal blk000004da_blk000004db_sig00001536 : STD_LOGIC; 
  signal blk000004da_blk000004db_sig00001535 : STD_LOGIC; 
  signal blk000004da_blk000004db_sig00001534 : STD_LOGIC; 
  signal blk000004da_blk000004db_sig00001533 : STD_LOGIC; 
  signal blk000004da_blk000004db_sig00001532 : STD_LOGIC; 
  signal blk000004da_blk000004db_sig00001531 : STD_LOGIC; 
  signal blk000004da_blk000004db_sig00001530 : STD_LOGIC; 
  signal blk000004da_blk000004db_sig0000152f : STD_LOGIC; 
  signal blk000004da_blk000004db_sig0000152e : STD_LOGIC; 
  signal blk000004da_blk000004db_sig0000152d : STD_LOGIC; 
  signal blk000004fa_blk000004fb_sig00001589 : STD_LOGIC; 
  signal blk000004fa_blk000004fb_sig00001588 : STD_LOGIC; 
  signal blk000004fa_blk000004fb_sig00001587 : STD_LOGIC; 
  signal blk000004fa_blk000004fb_sig00001586 : STD_LOGIC; 
  signal blk000004fa_blk000004fb_sig00001585 : STD_LOGIC; 
  signal blk000004fa_blk000004fb_sig00001584 : STD_LOGIC; 
  signal blk000004fa_blk000004fb_sig00001583 : STD_LOGIC; 
  signal blk000004fa_blk000004fb_sig00001582 : STD_LOGIC; 
  signal blk000004fa_blk000004fb_sig00001581 : STD_LOGIC; 
  signal blk000004fa_blk000004fb_sig00001580 : STD_LOGIC; 
  signal blk000004fa_blk000004fb_sig0000157f : STD_LOGIC; 
  signal blk000004fa_blk000004fb_sig0000157e : STD_LOGIC; 
  signal blk000004fa_blk000004fb_sig0000157d : STD_LOGIC; 
  signal blk000004fa_blk000004fb_sig0000157c : STD_LOGIC; 
  signal blk000004fa_blk000004fb_sig0000157b : STD_LOGIC; 
  signal blk000004fa_blk000004fb_sig0000157a : STD_LOGIC; 
  signal blk0000051a_blk0000051b_sig000015d6 : STD_LOGIC; 
  signal blk0000051a_blk0000051b_sig000015d5 : STD_LOGIC; 
  signal blk0000051a_blk0000051b_sig000015d4 : STD_LOGIC; 
  signal blk0000051a_blk0000051b_sig000015d3 : STD_LOGIC; 
  signal blk0000051a_blk0000051b_sig000015d2 : STD_LOGIC; 
  signal blk0000051a_blk0000051b_sig000015d1 : STD_LOGIC; 
  signal blk0000051a_blk0000051b_sig000015d0 : STD_LOGIC; 
  signal blk0000051a_blk0000051b_sig000015cf : STD_LOGIC; 
  signal blk0000051a_blk0000051b_sig000015ce : STD_LOGIC; 
  signal blk0000051a_blk0000051b_sig000015cd : STD_LOGIC; 
  signal blk0000051a_blk0000051b_sig000015cc : STD_LOGIC; 
  signal blk0000051a_blk0000051b_sig000015cb : STD_LOGIC; 
  signal blk0000051a_blk0000051b_sig000015ca : STD_LOGIC; 
  signal blk0000051a_blk0000051b_sig000015c9 : STD_LOGIC; 
  signal blk0000051a_blk0000051b_sig000015c8 : STD_LOGIC; 
  signal blk0000051a_blk0000051b_sig000015c7 : STD_LOGIC; 
  signal blk0000053a_sig0000162c : STD_LOGIC; 
  signal blk0000053a_sig0000162b : STD_LOGIC; 
  signal blk0000053a_sig0000162a : STD_LOGIC; 
  signal blk0000053a_sig00001629 : STD_LOGIC; 
  signal blk0000053a_sig00001628 : STD_LOGIC; 
  signal blk0000053a_sig00001627 : STD_LOGIC; 
  signal blk0000053a_sig00001626 : STD_LOGIC; 
  signal blk0000053a_sig00001625 : STD_LOGIC; 
  signal blk0000053a_sig00001624 : STD_LOGIC; 
  signal blk0000053a_sig00001623 : STD_LOGIC; 
  signal blk0000053a_sig00001622 : STD_LOGIC; 
  signal blk0000053a_sig00001621 : STD_LOGIC; 
  signal blk0000053a_sig00001620 : STD_LOGIC; 
  signal blk0000053a_sig0000161f : STD_LOGIC; 
  signal blk0000053a_sig0000161e : STD_LOGIC; 
  signal blk0000053a_sig0000161d : STD_LOGIC; 
  signal blk0000053a_sig0000161c : STD_LOGIC; 
  signal blk0000053a_sig0000161b : STD_LOGIC; 
  signal blk0000053a_sig0000161a : STD_LOGIC; 
  signal blk0000053a_sig00001619 : STD_LOGIC; 
  signal blk0000053a_sig00001618 : STD_LOGIC; 
  signal blk0000053a_sig00001617 : STD_LOGIC; 
  signal blk0000053a_sig00001616 : STD_LOGIC; 
  signal blk0000053a_sig00001615 : STD_LOGIC; 
  signal blk0000053a_sig00001614 : STD_LOGIC; 
  signal blk0000053a_sig00001613 : STD_LOGIC; 
  signal blk0000053a_sig00001612 : STD_LOGIC; 
  signal blk0000053a_sig00001611 : STD_LOGIC; 
  signal blk0000053a_sig00001610 : STD_LOGIC; 
  signal blk0000053a_sig0000160f : STD_LOGIC; 
  signal blk0000053a_sig0000160e : STD_LOGIC; 
  signal blk0000053a_sig0000160d : STD_LOGIC; 
  signal blk0000053a_sig0000160c : STD_LOGIC; 
  signal blk0000053a_sig0000160b : STD_LOGIC; 
  signal blk0000053a_sig0000160a : STD_LOGIC; 
  signal blk0000053a_sig00001609 : STD_LOGIC; 
  signal blk0000053a_sig00001608 : STD_LOGIC; 
  signal blk0000053a_sig00001607 : STD_LOGIC; 
  signal blk0000053a_sig00001606 : STD_LOGIC; 
  signal blk0000053a_sig00001605 : STD_LOGIC; 
  signal blk0000053a_sig00001604 : STD_LOGIC; 
  signal blk0000053a_sig00001603 : STD_LOGIC; 
  signal blk00000573_sig00001682 : STD_LOGIC; 
  signal blk00000573_sig00001681 : STD_LOGIC; 
  signal blk00000573_sig00001680 : STD_LOGIC; 
  signal blk00000573_sig0000167f : STD_LOGIC; 
  signal blk00000573_sig0000167e : STD_LOGIC; 
  signal blk00000573_sig0000167d : STD_LOGIC; 
  signal blk00000573_sig0000167c : STD_LOGIC; 
  signal blk00000573_sig0000167b : STD_LOGIC; 
  signal blk00000573_sig0000167a : STD_LOGIC; 
  signal blk00000573_sig00001679 : STD_LOGIC; 
  signal blk00000573_sig00001678 : STD_LOGIC; 
  signal blk00000573_sig00001677 : STD_LOGIC; 
  signal blk00000573_sig00001676 : STD_LOGIC; 
  signal blk00000573_sig00001675 : STD_LOGIC; 
  signal blk00000573_sig00001674 : STD_LOGIC; 
  signal blk00000573_sig00001673 : STD_LOGIC; 
  signal blk00000573_sig00001672 : STD_LOGIC; 
  signal blk00000573_sig00001671 : STD_LOGIC; 
  signal blk00000573_sig00001670 : STD_LOGIC; 
  signal blk00000573_sig0000166f : STD_LOGIC; 
  signal blk00000573_sig0000166e : STD_LOGIC; 
  signal blk00000573_sig0000166d : STD_LOGIC; 
  signal blk00000573_sig0000166c : STD_LOGIC; 
  signal blk00000573_sig0000166b : STD_LOGIC; 
  signal blk00000573_sig0000166a : STD_LOGIC; 
  signal blk00000573_sig00001669 : STD_LOGIC; 
  signal blk00000573_sig00001668 : STD_LOGIC; 
  signal blk00000573_sig00001667 : STD_LOGIC; 
  signal blk00000573_sig00001666 : STD_LOGIC; 
  signal blk00000573_sig00001665 : STD_LOGIC; 
  signal blk00000573_sig00001664 : STD_LOGIC; 
  signal blk00000573_sig00001663 : STD_LOGIC; 
  signal blk00000573_sig00001662 : STD_LOGIC; 
  signal blk00000573_sig00001661 : STD_LOGIC; 
  signal blk00000573_sig00001660 : STD_LOGIC; 
  signal blk00000573_sig0000165f : STD_LOGIC; 
  signal blk00000573_sig0000165e : STD_LOGIC; 
  signal blk00000573_sig0000165d : STD_LOGIC; 
  signal blk00000573_sig0000165c : STD_LOGIC; 
  signal blk00000573_sig0000165b : STD_LOGIC; 
  signal blk00000573_sig0000165a : STD_LOGIC; 
  signal blk00000573_sig00001659 : STD_LOGIC; 
  signal blk000005ac_blk000005ad_sig000016a6 : STD_LOGIC; 
  signal blk000005ac_blk000005ad_sig000016a5 : STD_LOGIC; 
  signal blk000005ac_blk000005ad_sig000016a4 : STD_LOGIC; 
  signal blk000005ac_blk000005ad_sig000016a3 : STD_LOGIC; 
  signal blk000005ac_blk000005ad_sig000016a2 : STD_LOGIC; 
  signal blk000005ac_blk000005ad_sig000016a1 : STD_LOGIC; 
  signal blk000005ac_blk000005ad_sig000016a0 : STD_LOGIC; 
  signal blk000005ac_blk000005ad_sig0000169f : STD_LOGIC; 
  signal blk000005bc_blk000005bd_sig000016b1 : STD_LOGIC; 
  signal blk000005bc_blk000005bd_sig000016b0 : STD_LOGIC; 
  signal blk000005bc_blk000005bd_sig000016af : STD_LOGIC; 
  signal blk000005c2_blk000005c3_sig000016c2 : STD_LOGIC; 
  signal blk000005c2_blk000005c3_sig000016c1 : STD_LOGIC; 
  signal blk000005cd_sig000016e4 : STD_LOGIC; 
  signal blk000005cd_sig000016e3 : STD_LOGIC; 
  signal blk000005cd_sig000016e2 : STD_LOGIC; 
  signal blk000005cd_sig000016e1 : STD_LOGIC; 
  signal blk000005cd_sig000016e0 : STD_LOGIC; 
  signal blk000005cd_sig000016df : STD_LOGIC; 
  signal blk000005cd_sig000016de : STD_LOGIC; 
  signal blk000005cd_sig000016dd : STD_LOGIC; 
  signal blk000005cd_sig000016dc : STD_LOGIC; 
  signal blk000005cd_sig000016db : STD_LOGIC; 
  signal blk000005cd_sig000016da : STD_LOGIC; 
  signal blk000005cd_sig000016d9 : STD_LOGIC; 
  signal blk000005cd_sig000016d8 : STD_LOGIC; 
  signal blk000005cd_sig000016d7 : STD_LOGIC; 
  signal blk000005cd_sig000016d6 : STD_LOGIC; 
  signal blk000005cd_sig000016d5 : STD_LOGIC; 
  signal blk000005cd_sig000016d4 : STD_LOGIC; 
  signal blk000005f1_sig0000174f : STD_LOGIC; 
  signal blk000005f1_sig0000174e : STD_LOGIC; 
  signal blk000005f1_sig0000174d : STD_LOGIC; 
  signal blk000005f1_sig0000174c : STD_LOGIC; 
  signal blk000005f1_sig0000174b : STD_LOGIC; 
  signal blk000005f1_sig0000174a : STD_LOGIC; 
  signal blk000005f1_sig00001749 : STD_LOGIC; 
  signal blk000005f1_sig00001748 : STD_LOGIC; 
  signal blk000005f1_sig00001747 : STD_LOGIC; 
  signal blk000005f1_sig00001746 : STD_LOGIC; 
  signal blk000005f1_sig00001745 : STD_LOGIC; 
  signal blk000005f1_sig00001744 : STD_LOGIC; 
  signal blk000005f1_sig00001743 : STD_LOGIC; 
  signal blk000005f1_sig00001742 : STD_LOGIC; 
  signal blk000005f1_sig00001741 : STD_LOGIC; 
  signal blk000005f1_sig00001740 : STD_LOGIC; 
  signal blk000005f1_sig0000173f : STD_LOGIC; 
  signal blk000005f1_sig0000173e : STD_LOGIC; 
  signal blk000005f1_sig0000173d : STD_LOGIC; 
  signal blk000005f1_sig0000173c : STD_LOGIC; 
  signal blk000005f1_sig0000173b : STD_LOGIC; 
  signal blk000005f1_sig0000173a : STD_LOGIC; 
  signal blk000005f1_sig00001739 : STD_LOGIC; 
  signal blk000005f1_sig00001738 : STD_LOGIC; 
  signal blk000005f1_sig00001737 : STD_LOGIC; 
  signal blk000005f1_sig00001736 : STD_LOGIC; 
  signal blk000005f1_sig00001735 : STD_LOGIC; 
  signal blk000005f1_sig00001734 : STD_LOGIC; 
  signal blk000005f1_sig00001733 : STD_LOGIC; 
  signal blk000005f1_sig00001732 : STD_LOGIC; 
  signal blk000005f1_sig00001731 : STD_LOGIC; 
  signal blk000005f1_sig00001730 : STD_LOGIC; 
  signal blk000005f1_sig0000172f : STD_LOGIC; 
  signal blk000005f1_sig0000172e : STD_LOGIC; 
  signal blk000005f1_sig0000172d : STD_LOGIC; 
  signal blk000005f1_sig0000172c : STD_LOGIC; 
  signal blk000005f1_sig0000172b : STD_LOGIC; 
  signal blk000005f1_sig0000172a : STD_LOGIC; 
  signal blk000005f1_sig00001729 : STD_LOGIC; 
  signal blk000005f1_sig00001728 : STD_LOGIC; 
  signal blk000005f1_sig00001727 : STD_LOGIC; 
  signal blk000005f1_sig00001726 : STD_LOGIC; 
  signal blk000005f1_sig00001725 : STD_LOGIC; 
  signal blk000005f1_sig00001724 : STD_LOGIC; 
  signal blk000005f1_sig00001723 : STD_LOGIC; 
  signal blk000005f1_sig00001722 : STD_LOGIC; 
  signal blk000005f1_sig00001721 : STD_LOGIC; 
  signal blk000005f1_sig00001720 : STD_LOGIC; 
  signal blk000005f1_sig0000171f : STD_LOGIC; 
  signal blk000005f1_sig0000171e : STD_LOGIC; 
  signal blk000005f1_sig0000171d : STD_LOGIC; 
  signal blk000005f1_sig0000171c : STD_LOGIC; 
  signal blk000005f1_sig0000171b : STD_LOGIC; 
  signal blk000005f1_sig0000171a : STD_LOGIC; 
  signal blk000005f1_sig00001719 : STD_LOGIC; 
  signal blk000005f1_sig00001718 : STD_LOGIC; 
  signal blk000005f1_sig00001717 : STD_LOGIC; 
  signal blk000005f1_sig00001716 : STD_LOGIC; 
  signal blk000005f1_sig00001715 : STD_LOGIC; 
  signal blk000005f1_sig00001714 : STD_LOGIC; 
  signal blk000005f1_sig000016f9 : STD_LOGIC; 
  signal blk000005f1_sig000016f8 : STD_LOGIC; 
  signal blk000005f1_sig000016f7 : STD_LOGIC; 
  signal blk000005f1_sig000016f6 : STD_LOGIC; 
  signal blk000005f1_sig000016f5 : STD_LOGIC; 
  signal blk000005f1_sig000016f4 : STD_LOGIC; 
  signal blk000005f1_sig000016f3 : STD_LOGIC; 
  signal blk000005f1_sig000016f2 : STD_LOGIC; 
  signal blk000005f1_sig000016f1 : STD_LOGIC; 
  signal blk000005f1_sig000016f0 : STD_LOGIC; 
  signal blk000005f1_sig000016ef : STD_LOGIC; 
  signal blk000005f1_sig000016ee : STD_LOGIC; 
  signal blk000005f1_sig000016ed : STD_LOGIC; 
  signal blk0000091a_blk0000091b_sig0000195f : STD_LOGIC; 
  signal blk0000091a_blk0000091b_sig0000195e : STD_LOGIC; 
  signal blk0000091a_blk0000091b_sig0000195d : STD_LOGIC; 
  signal blk0000092d_sig0000197f : STD_LOGIC; 
  signal blk0000092d_sig0000197e : STD_LOGIC; 
  signal blk0000092d_sig0000197d : STD_LOGIC; 
  signal blk0000092d_sig0000197c : STD_LOGIC; 
  signal blk0000092d_sig0000197b : STD_LOGIC; 
  signal blk0000092d_sig0000197a : STD_LOGIC; 
  signal blk0000092d_sig00001979 : STD_LOGIC; 
  signal blk0000092d_sig00001978 : STD_LOGIC; 
  signal blk0000092d_sig00001977 : STD_LOGIC; 
  signal blk0000092d_sig00001976 : STD_LOGIC; 
  signal blk0000092d_sig00001975 : STD_LOGIC; 
  signal blk0000092d_sig00001974 : STD_LOGIC; 
  signal blk0000092d_sig00001973 : STD_LOGIC; 
  signal blk0000092d_sig00001972 : STD_LOGIC; 
  signal blk0000092d_sig00001971 : STD_LOGIC; 
  signal blk0000092d_sig00001970 : STD_LOGIC; 
  signal blk00000955_sig0000199f : STD_LOGIC; 
  signal blk00000955_sig0000199e : STD_LOGIC; 
  signal blk00000955_sig0000199d : STD_LOGIC; 
  signal blk00000955_sig0000199c : STD_LOGIC; 
  signal blk00000955_sig0000199b : STD_LOGIC; 
  signal blk00000955_sig0000199a : STD_LOGIC; 
  signal blk00000955_sig00001999 : STD_LOGIC; 
  signal blk00000955_sig00001998 : STD_LOGIC; 
  signal blk00000955_sig00001997 : STD_LOGIC; 
  signal blk00000955_sig00001996 : STD_LOGIC; 
  signal blk00000955_sig00001995 : STD_LOGIC; 
  signal blk00000955_sig00001994 : STD_LOGIC; 
  signal blk00000955_sig00001993 : STD_LOGIC; 
  signal blk00000955_sig00001992 : STD_LOGIC; 
  signal blk00000955_sig00001991 : STD_LOGIC; 
  signal blk00000955_sig00001990 : STD_LOGIC; 
  signal blk000009b1_blk000009b2_sig000019e2 : STD_LOGIC; 
  signal blk000009b1_blk000009b2_sig000019e1 : STD_LOGIC; 
  signal blk000009b1_blk000009b2_sig000019e0 : STD_LOGIC; 
  signal blk000009b1_blk000009b2_sig000019df : STD_LOGIC; 
  signal blk000009b1_blk000009b2_sig000019de : STD_LOGIC; 
  signal blk000009b1_blk000009b2_sig000019dd : STD_LOGIC; 
  signal blk000009b1_blk000009b2_sig000019dc : STD_LOGIC; 
  signal blk000009b1_blk000009b2_sig000019db : STD_LOGIC; 
  signal blk000009b1_blk000009b2_sig000019da : STD_LOGIC; 
  signal blk000009b1_blk000009b2_sig000019d9 : STD_LOGIC; 
  signal blk000009b1_blk000009b2_sig000019d8 : STD_LOGIC; 
  signal blk000009b1_blk000009b2_sig000019d7 : STD_LOGIC; 
  signal blk000009b1_blk000009b2_sig000019d6 : STD_LOGIC; 
  signal blk000009b1_blk000009b2_sig000019d5 : STD_LOGIC; 
  signal blk000009cd_blk000009ce_sig00001a25 : STD_LOGIC; 
  signal blk000009cd_blk000009ce_sig00001a24 : STD_LOGIC; 
  signal blk000009cd_blk000009ce_sig00001a23 : STD_LOGIC; 
  signal blk000009cd_blk000009ce_sig00001a22 : STD_LOGIC; 
  signal blk000009cd_blk000009ce_sig00001a21 : STD_LOGIC; 
  signal blk000009cd_blk000009ce_sig00001a20 : STD_LOGIC; 
  signal blk000009cd_blk000009ce_sig00001a1f : STD_LOGIC; 
  signal blk000009cd_blk000009ce_sig00001a1e : STD_LOGIC; 
  signal blk000009cd_blk000009ce_sig00001a1d : STD_LOGIC; 
  signal blk000009cd_blk000009ce_sig00001a1c : STD_LOGIC; 
  signal blk000009cd_blk000009ce_sig00001a1b : STD_LOGIC; 
  signal blk000009cd_blk000009ce_sig00001a1a : STD_LOGIC; 
  signal blk000009cd_blk000009ce_sig00001a19 : STD_LOGIC; 
  signal blk000009cd_blk000009ce_sig00001a18 : STD_LOGIC; 
  signal blk000009e9_blk000009ea_sig00001a30 : STD_LOGIC; 
  signal blk000009e9_blk000009ea_sig00001a2f : STD_LOGIC; 
  signal blk000009e9_blk000009ea_sig00001a2e : STD_LOGIC; 
  signal blk000009ef_sig00001a7e : STD_LOGIC; 
  signal blk000009ef_sig00001a7d : STD_LOGIC; 
  signal blk000009ef_sig00001a7c : STD_LOGIC; 
  signal blk000009ef_sig00001a7b : STD_LOGIC; 
  signal blk000009ef_sig00001a7a : STD_LOGIC; 
  signal blk000009ef_sig00001a79 : STD_LOGIC; 
  signal blk000009ef_sig00001a78 : STD_LOGIC; 
  signal blk000009ef_sig00001a77 : STD_LOGIC; 
  signal blk000009ef_sig00001a76 : STD_LOGIC; 
  signal blk000009ef_sig00001a75 : STD_LOGIC; 
  signal blk000009ef_sig00001a74 : STD_LOGIC; 
  signal blk000009ef_sig00001a73 : STD_LOGIC; 
  signal blk000009ef_sig00001a72 : STD_LOGIC; 
  signal blk000009ef_sig00001a71 : STD_LOGIC; 
  signal blk000009ef_sig00001a70 : STD_LOGIC; 
  signal blk000009ef_sig00001a6f : STD_LOGIC; 
  signal blk000009ef_sig00001a6e : STD_LOGIC; 
  signal blk000009ef_sig00001a6d : STD_LOGIC; 
  signal blk000009ef_sig00001a6c : STD_LOGIC; 
  signal blk000009ef_sig00001a6b : STD_LOGIC; 
  signal blk000009ef_sig00001a6a : STD_LOGIC; 
  signal blk000009ef_sig00001a69 : STD_LOGIC; 
  signal blk000009ef_sig00001a68 : STD_LOGIC; 
  signal blk000009ef_sig00001a67 : STD_LOGIC; 
  signal blk000009ef_sig00001a66 : STD_LOGIC; 
  signal blk000009ef_sig00001a65 : STD_LOGIC; 
  signal blk000009ef_sig00001a64 : STD_LOGIC; 
  signal blk000009ef_sig00001a63 : STD_LOGIC; 
  signal blk000009ef_sig00001a62 : STD_LOGIC; 
  signal blk000009ef_sig00001a61 : STD_LOGIC; 
  signal blk000009ef_sig00001a60 : STD_LOGIC; 
  signal blk000009ef_sig00001a5f : STD_LOGIC; 
  signal blk000009ef_sig00001a5e : STD_LOGIC; 
  signal blk000009ef_sig00001a5d : STD_LOGIC; 
  signal blk000009ef_sig00001a5c : STD_LOGIC; 
  signal blk000009ef_sig00001a5b : STD_LOGIC; 
  signal blk000009ef_sig00001a5a : STD_LOGIC; 
  signal blk000009ef_sig00001a59 : STD_LOGIC; 
  signal blk000009ef_sig00001a58 : STD_LOGIC; 
  signal blk00000a24_sig00001acc : STD_LOGIC; 
  signal blk00000a24_sig00001acb : STD_LOGIC; 
  signal blk00000a24_sig00001aca : STD_LOGIC; 
  signal blk00000a24_sig00001ac9 : STD_LOGIC; 
  signal blk00000a24_sig00001ac8 : STD_LOGIC; 
  signal blk00000a24_sig00001ac7 : STD_LOGIC; 
  signal blk00000a24_sig00001ac6 : STD_LOGIC; 
  signal blk00000a24_sig00001ac5 : STD_LOGIC; 
  signal blk00000a24_sig00001ac4 : STD_LOGIC; 
  signal blk00000a24_sig00001ac3 : STD_LOGIC; 
  signal blk00000a24_sig00001ac2 : STD_LOGIC; 
  signal blk00000a24_sig00001ac1 : STD_LOGIC; 
  signal blk00000a24_sig00001ac0 : STD_LOGIC; 
  signal blk00000a24_sig00001abf : STD_LOGIC; 
  signal blk00000a24_sig00001abe : STD_LOGIC; 
  signal blk00000a24_sig00001abd : STD_LOGIC; 
  signal blk00000a24_sig00001abc : STD_LOGIC; 
  signal blk00000a24_sig00001abb : STD_LOGIC; 
  signal blk00000a24_sig00001aba : STD_LOGIC; 
  signal blk00000a24_sig00001ab9 : STD_LOGIC; 
  signal blk00000a24_sig00001ab8 : STD_LOGIC; 
  signal blk00000a24_sig00001ab7 : STD_LOGIC; 
  signal blk00000a24_sig00001ab6 : STD_LOGIC; 
  signal blk00000a24_sig00001ab5 : STD_LOGIC; 
  signal blk00000a24_sig00001ab4 : STD_LOGIC; 
  signal blk00000a24_sig00001ab3 : STD_LOGIC; 
  signal blk00000a24_sig00001ab2 : STD_LOGIC; 
  signal blk00000a24_sig00001ab1 : STD_LOGIC; 
  signal blk00000a24_sig00001ab0 : STD_LOGIC; 
  signal blk00000a24_sig00001aaf : STD_LOGIC; 
  signal blk00000a24_sig00001aae : STD_LOGIC; 
  signal blk00000a24_sig00001aad : STD_LOGIC; 
  signal blk00000a24_sig00001aac : STD_LOGIC; 
  signal blk00000a24_sig00001aab : STD_LOGIC; 
  signal blk00000a24_sig00001aaa : STD_LOGIC; 
  signal blk00000a24_sig00001aa9 : STD_LOGIC; 
  signal blk00000a24_sig00001aa8 : STD_LOGIC; 
  signal blk00000a24_sig00001aa7 : STD_LOGIC; 
  signal blk00000a24_sig00001aa6 : STD_LOGIC; 
  signal blk00000a59_blk00000a5a_sig00001b14 : STD_LOGIC; 
  signal blk00000a59_blk00000a5a_sig00001b13 : STD_LOGIC; 
  signal blk00000a59_blk00000a5a_sig00001b12 : STD_LOGIC; 
  signal blk00000a59_blk00000a5a_sig00001b11 : STD_LOGIC; 
  signal blk00000a59_blk00000a5a_sig00001b10 : STD_LOGIC; 
  signal blk00000a59_blk00000a5a_sig00001b0f : STD_LOGIC; 
  signal blk00000a59_blk00000a5a_sig00001b0e : STD_LOGIC; 
  signal blk00000a59_blk00000a5a_sig00001b0d : STD_LOGIC; 
  signal blk00000a59_blk00000a5a_sig00001b0c : STD_LOGIC; 
  signal blk00000a59_blk00000a5a_sig00001b0b : STD_LOGIC; 
  signal blk00000a59_blk00000a5a_sig00001b0a : STD_LOGIC; 
  signal blk00000a59_blk00000a5a_sig00001b09 : STD_LOGIC; 
  signal blk00000a59_blk00000a5a_sig00001b08 : STD_LOGIC; 
  signal blk00000a59_blk00000a5a_sig00001b07 : STD_LOGIC; 
  signal blk00000a59_blk00000a5a_sig00001b06 : STD_LOGIC; 
  signal blk00000a77_blk00000a78_sig00001b5c : STD_LOGIC; 
  signal blk00000a77_blk00000a78_sig00001b5b : STD_LOGIC; 
  signal blk00000a77_blk00000a78_sig00001b5a : STD_LOGIC; 
  signal blk00000a77_blk00000a78_sig00001b59 : STD_LOGIC; 
  signal blk00000a77_blk00000a78_sig00001b58 : STD_LOGIC; 
  signal blk00000a77_blk00000a78_sig00001b57 : STD_LOGIC; 
  signal blk00000a77_blk00000a78_sig00001b56 : STD_LOGIC; 
  signal blk00000a77_blk00000a78_sig00001b55 : STD_LOGIC; 
  signal blk00000a77_blk00000a78_sig00001b54 : STD_LOGIC; 
  signal blk00000a77_blk00000a78_sig00001b53 : STD_LOGIC; 
  signal blk00000a77_blk00000a78_sig00001b52 : STD_LOGIC; 
  signal blk00000a77_blk00000a78_sig00001b51 : STD_LOGIC; 
  signal blk00000a77_blk00000a78_sig00001b50 : STD_LOGIC; 
  signal blk00000a77_blk00000a78_sig00001b4f : STD_LOGIC; 
  signal blk00000a77_blk00000a78_sig00001b4e : STD_LOGIC; 
  signal blk00000a95_sig00001b64 : STD_LOGIC; 
  signal blk00000a95_sig00001b63 : STD_LOGIC; 
  signal blk00000a95_blk00000a96_sig00001b70 : STD_LOGIC; 
  signal blk00000a95_blk00000a96_sig00001b6f : STD_LOGIC; 
  signal blk00000a95_blk00000a96_sig00001b6e : STD_LOGIC; 
  signal blk00000a95_blk00000a96_sig00001b6d : STD_LOGIC; 
  signal blk00000a9d_blk00000a9e_sig00001b7b : STD_LOGIC; 
  signal blk00000a9d_blk00000a9e_sig00001b7a : STD_LOGIC; 
  signal blk00000a9d_blk00000a9e_sig00001b79 : STD_LOGIC; 
  signal blk00000aa3_blk00000aa4_sig00001b86 : STD_LOGIC; 
  signal blk00000aa3_blk00000aa4_sig00001b85 : STD_LOGIC; 
  signal blk00000aa3_blk00000aa4_sig00001b84 : STD_LOGIC; 
  signal blk00000aa9_blk00000aaa_sig00001b91 : STD_LOGIC; 
  signal blk00000aa9_blk00000aaa_sig00001b90 : STD_LOGIC; 
  signal blk00000aa9_blk00000aaa_sig00001b8f : STD_LOGIC; 
  signal blk00000aaf_blk00000ab0_sig00001ba1 : STD_LOGIC; 
  signal blk00000aaf_blk00000ab0_sig00001ba0 : STD_LOGIC; 
  signal blk00000aaf_blk00000ab0_sig00001b9f : STD_LOGIC; 
  signal blk00000aaf_blk00000ab0_sig00001b9e : STD_LOGIC; 
  signal blk00000ab7_blk00000ab8_sig00001bb1 : STD_LOGIC; 
  signal blk00000ab7_blk00000ab8_sig00001bb0 : STD_LOGIC; 
  signal blk00000ab7_blk00000ab8_sig00001baf : STD_LOGIC; 
  signal blk00000ab7_blk00000ab8_sig00001bae : STD_LOGIC; 
  signal blk00000abf_blk00000ac0_sig00001bd5 : STD_LOGIC; 
  signal blk00000abf_blk00000ac0_sig00001bd4 : STD_LOGIC; 
  signal blk00000abf_blk00000ac0_sig00001bd3 : STD_LOGIC; 
  signal blk00000abf_blk00000ac0_sig00001bd2 : STD_LOGIC; 
  signal blk00000abf_blk00000ac0_sig00001bd1 : STD_LOGIC; 
  signal blk00000abf_blk00000ac0_sig00001bd0 : STD_LOGIC; 
  signal blk00000abf_blk00000ac0_sig00001bcf : STD_LOGIC; 
  signal blk00000abf_blk00000ac0_sig00001bce : STD_LOGIC; 
  signal blk00000acf_sig00001bdf : STD_LOGIC; 
  signal blk00000acf_sig00001bde : STD_LOGIC; 
  signal blk00000acf_blk00000ad0_sig00001be9 : STD_LOGIC; 
  signal blk00000acf_blk00000ad0_sig00001be8 : STD_LOGIC; 
  signal blk00000acf_blk00000ad0_sig00001be7 : STD_LOGIC; 
  signal blk00000acf_blk00000ad0_sig00001be6 : STD_LOGIC; 
  signal blk00000ad7_sig00001c3f : STD_LOGIC; 
  signal blk00000ad7_sig00001c3e : STD_LOGIC; 
  signal blk00000ad7_sig00001c3d : STD_LOGIC; 
  signal blk00000ad7_sig00001c3c : STD_LOGIC; 
  signal blk00000ad7_sig00001c3b : STD_LOGIC; 
  signal blk00000ad7_sig00001c3a : STD_LOGIC; 
  signal blk00000ad7_sig00001c39 : STD_LOGIC; 
  signal blk00000ad7_sig00001c38 : STD_LOGIC; 
  signal blk00000ad7_sig00001c37 : STD_LOGIC; 
  signal blk00000ad7_sig00001c36 : STD_LOGIC; 
  signal blk00000ad7_sig00001c35 : STD_LOGIC; 
  signal blk00000ad7_sig00001c34 : STD_LOGIC; 
  signal blk00000ad7_sig00001c33 : STD_LOGIC; 
  signal blk00000ad7_sig00001c32 : STD_LOGIC; 
  signal blk00000ad7_sig00001c31 : STD_LOGIC; 
  signal blk00000ad7_sig00001c30 : STD_LOGIC; 
  signal blk00000ad7_sig00001c2f : STD_LOGIC; 
  signal blk00000ad7_sig00001c2e : STD_LOGIC; 
  signal blk00000ad7_sig00001c2d : STD_LOGIC; 
  signal blk00000ad7_sig00001c2c : STD_LOGIC; 
  signal blk00000ad7_sig00001c2b : STD_LOGIC; 
  signal blk00000ad7_sig00001c2a : STD_LOGIC; 
  signal blk00000ad7_sig00001c29 : STD_LOGIC; 
  signal blk00000ad7_sig00001c28 : STD_LOGIC; 
  signal blk00000ad7_sig00001c27 : STD_LOGIC; 
  signal blk00000ad7_sig00001c26 : STD_LOGIC; 
  signal blk00000ad7_sig00001c25 : STD_LOGIC; 
  signal blk00000ad7_sig00001c24 : STD_LOGIC; 
  signal blk00000ad7_sig00001c23 : STD_LOGIC; 
  signal blk00000ad7_sig00001c22 : STD_LOGIC; 
  signal blk00000ad7_sig00001c21 : STD_LOGIC; 
  signal blk00000ad7_sig00001c20 : STD_LOGIC; 
  signal blk00000ad7_sig00001c1f : STD_LOGIC; 
  signal blk00000ad7_sig00001c1e : STD_LOGIC; 
  signal blk00000ad7_sig00001c1d : STD_LOGIC; 
  signal blk00000ad7_sig00001c1c : STD_LOGIC; 
  signal blk00000ad7_sig00001c1b : STD_LOGIC; 
  signal blk00000ad7_sig00001c1a : STD_LOGIC; 
  signal blk00000ad7_sig00001c19 : STD_LOGIC; 
  signal blk00000ad7_sig00001c18 : STD_LOGIC; 
  signal blk00000ad7_sig00001c17 : STD_LOGIC; 
  signal blk00000ad7_sig00001c16 : STD_LOGIC; 
  signal blk00000b10_sig00001c95 : STD_LOGIC; 
  signal blk00000b10_sig00001c94 : STD_LOGIC; 
  signal blk00000b10_sig00001c93 : STD_LOGIC; 
  signal blk00000b10_sig00001c92 : STD_LOGIC; 
  signal blk00000b10_sig00001c91 : STD_LOGIC; 
  signal blk00000b10_sig00001c90 : STD_LOGIC; 
  signal blk00000b10_sig00001c8f : STD_LOGIC; 
  signal blk00000b10_sig00001c8e : STD_LOGIC; 
  signal blk00000b10_sig00001c8d : STD_LOGIC; 
  signal blk00000b10_sig00001c8c : STD_LOGIC; 
  signal blk00000b10_sig00001c8b : STD_LOGIC; 
  signal blk00000b10_sig00001c8a : STD_LOGIC; 
  signal blk00000b10_sig00001c89 : STD_LOGIC; 
  signal blk00000b10_sig00001c88 : STD_LOGIC; 
  signal blk00000b10_sig00001c87 : STD_LOGIC; 
  signal blk00000b10_sig00001c86 : STD_LOGIC; 
  signal blk00000b10_sig00001c85 : STD_LOGIC; 
  signal blk00000b10_sig00001c84 : STD_LOGIC; 
  signal blk00000b10_sig00001c83 : STD_LOGIC; 
  signal blk00000b10_sig00001c82 : STD_LOGIC; 
  signal blk00000b10_sig00001c81 : STD_LOGIC; 
  signal blk00000b10_sig00001c80 : STD_LOGIC; 
  signal blk00000b10_sig00001c7f : STD_LOGIC; 
  signal blk00000b10_sig00001c7e : STD_LOGIC; 
  signal blk00000b10_sig00001c7d : STD_LOGIC; 
  signal blk00000b10_sig00001c7c : STD_LOGIC; 
  signal blk00000b10_sig00001c7b : STD_LOGIC; 
  signal blk00000b10_sig00001c7a : STD_LOGIC; 
  signal blk00000b10_sig00001c79 : STD_LOGIC; 
  signal blk00000b10_sig00001c78 : STD_LOGIC; 
  signal blk00000b10_sig00001c77 : STD_LOGIC; 
  signal blk00000b10_sig00001c76 : STD_LOGIC; 
  signal blk00000b10_sig00001c75 : STD_LOGIC; 
  signal blk00000b10_sig00001c74 : STD_LOGIC; 
  signal blk00000b10_sig00001c73 : STD_LOGIC; 
  signal blk00000b10_sig00001c72 : STD_LOGIC; 
  signal blk00000b10_sig00001c71 : STD_LOGIC; 
  signal blk00000b10_sig00001c70 : STD_LOGIC; 
  signal blk00000b10_sig00001c6f : STD_LOGIC; 
  signal blk00000b10_sig00001c6e : STD_LOGIC; 
  signal blk00000b10_sig00001c6d : STD_LOGIC; 
  signal blk00000b10_sig00001c6c : STD_LOGIC; 
  signal blk00000b49_blk00000b4a_sig00001ca6 : STD_LOGIC; 
  signal blk00000b49_blk00000b4a_sig00001ca5 : STD_LOGIC; 
  signal blk00000b4e_blk00000b4f_sig00001cb7 : STD_LOGIC; 
  signal blk00000b4e_blk00000b4f_sig00001cb6 : STD_LOGIC; 
  signal blk00000b53_blk00000b54_sig00001cc3 : STD_LOGIC; 
  signal blk00000b53_blk00000b54_sig00001cc2 : STD_LOGIC; 
  signal blk00000b53_blk00000b54_sig00001cc1 : STD_LOGIC; 
  signal blk00000c06_blk00000c07_sig00001d10 : STD_LOGIC; 
  signal blk00000c06_blk00000c07_sig00001d0f : STD_LOGIC; 
  signal blk00000c06_blk00000c07_sig00001d0e : STD_LOGIC; 
  signal blk00000c06_blk00000c07_sig00001d0d : STD_LOGIC; 
  signal blk00000c06_blk00000c07_sig00001d0c : STD_LOGIC; 
  signal blk00000c06_blk00000c07_sig00001d0b : STD_LOGIC; 
  signal blk00000c06_blk00000c07_sig00001d0a : STD_LOGIC; 
  signal blk00000c06_blk00000c07_sig00001d09 : STD_LOGIC; 
  signal blk00000c06_blk00000c07_sig00001d08 : STD_LOGIC; 
  signal blk00000c06_blk00000c07_sig00001d07 : STD_LOGIC; 
  signal blk00000c06_blk00000c07_sig00001d06 : STD_LOGIC; 
  signal blk00000c06_blk00000c07_sig00001d05 : STD_LOGIC; 
  signal blk00000c06_blk00000c07_sig00001d04 : STD_LOGIC; 
  signal blk00000c06_blk00000c07_sig00001d03 : STD_LOGIC; 
  signal blk00000c06_blk00000c07_sig00001d02 : STD_LOGIC; 
  signal blk00000c06_blk00000c07_sig00001d01 : STD_LOGIC; 
  signal blk00000c26_blk00000c27_sig00001d5d : STD_LOGIC; 
  signal blk00000c26_blk00000c27_sig00001d5c : STD_LOGIC; 
  signal blk00000c26_blk00000c27_sig00001d5b : STD_LOGIC; 
  signal blk00000c26_blk00000c27_sig00001d5a : STD_LOGIC; 
  signal blk00000c26_blk00000c27_sig00001d59 : STD_LOGIC; 
  signal blk00000c26_blk00000c27_sig00001d58 : STD_LOGIC; 
  signal blk00000c26_blk00000c27_sig00001d57 : STD_LOGIC; 
  signal blk00000c26_blk00000c27_sig00001d56 : STD_LOGIC; 
  signal blk00000c26_blk00000c27_sig00001d55 : STD_LOGIC; 
  signal blk00000c26_blk00000c27_sig00001d54 : STD_LOGIC; 
  signal blk00000c26_blk00000c27_sig00001d53 : STD_LOGIC; 
  signal blk00000c26_blk00000c27_sig00001d52 : STD_LOGIC; 
  signal blk00000c26_blk00000c27_sig00001d51 : STD_LOGIC; 
  signal blk00000c26_blk00000c27_sig00001d50 : STD_LOGIC; 
  signal blk00000c26_blk00000c27_sig00001d4f : STD_LOGIC; 
  signal blk00000c26_blk00000c27_sig00001d4e : STD_LOGIC; 
  signal blk00000c46_blk00000c47_sig00001daa : STD_LOGIC; 
  signal blk00000c46_blk00000c47_sig00001da9 : STD_LOGIC; 
  signal blk00000c46_blk00000c47_sig00001da8 : STD_LOGIC; 
  signal blk00000c46_blk00000c47_sig00001da7 : STD_LOGIC; 
  signal blk00000c46_blk00000c47_sig00001da6 : STD_LOGIC; 
  signal blk00000c46_blk00000c47_sig00001da5 : STD_LOGIC; 
  signal blk00000c46_blk00000c47_sig00001da4 : STD_LOGIC; 
  signal blk00000c46_blk00000c47_sig00001da3 : STD_LOGIC; 
  signal blk00000c46_blk00000c47_sig00001da2 : STD_LOGIC; 
  signal blk00000c46_blk00000c47_sig00001da1 : STD_LOGIC; 
  signal blk00000c46_blk00000c47_sig00001da0 : STD_LOGIC; 
  signal blk00000c46_blk00000c47_sig00001d9f : STD_LOGIC; 
  signal blk00000c46_blk00000c47_sig00001d9e : STD_LOGIC; 
  signal blk00000c46_blk00000c47_sig00001d9d : STD_LOGIC; 
  signal blk00000c46_blk00000c47_sig00001d9c : STD_LOGIC; 
  signal blk00000c46_blk00000c47_sig00001d9b : STD_LOGIC; 
  signal blk00000c66_blk00000c67_sig00001df7 : STD_LOGIC; 
  signal blk00000c66_blk00000c67_sig00001df6 : STD_LOGIC; 
  signal blk00000c66_blk00000c67_sig00001df5 : STD_LOGIC; 
  signal blk00000c66_blk00000c67_sig00001df4 : STD_LOGIC; 
  signal blk00000c66_blk00000c67_sig00001df3 : STD_LOGIC; 
  signal blk00000c66_blk00000c67_sig00001df2 : STD_LOGIC; 
  signal blk00000c66_blk00000c67_sig00001df1 : STD_LOGIC; 
  signal blk00000c66_blk00000c67_sig00001df0 : STD_LOGIC; 
  signal blk00000c66_blk00000c67_sig00001def : STD_LOGIC; 
  signal blk00000c66_blk00000c67_sig00001dee : STD_LOGIC; 
  signal blk00000c66_blk00000c67_sig00001ded : STD_LOGIC; 
  signal blk00000c66_blk00000c67_sig00001dec : STD_LOGIC; 
  signal blk00000c66_blk00000c67_sig00001deb : STD_LOGIC; 
  signal blk00000c66_blk00000c67_sig00001dea : STD_LOGIC; 
  signal blk00000c66_blk00000c67_sig00001de9 : STD_LOGIC; 
  signal blk00000c66_blk00000c67_sig00001de8 : STD_LOGIC; 
  signal blk00000c86_blk00000c87_sig00001e11 : STD_LOGIC; 
  signal blk00000c86_blk00000c87_sig00001e10 : STD_LOGIC; 
  signal blk00000c86_blk00000c87_sig00001e0f : STD_LOGIC; 
  signal blk00000c86_blk00000c87_sig00001e0e : STD_LOGIC; 
  signal blk00000c86_blk00000c87_sig00001e0d : STD_LOGIC; 
  signal blk00000c86_blk00000c87_sig00001e0c : STD_LOGIC; 
  signal blk00000c92_blk00000c93_sig00001e22 : STD_LOGIC; 
  signal blk00000c92_blk00000c93_sig00001e21 : STD_LOGIC; 
  signal blk00000c9b_sig00001e38 : STD_LOGIC; 
  signal blk00000c9b_sig00001e37 : STD_LOGIC; 
  signal blk00000c9b_sig00001e36 : STD_LOGIC; 
  signal blk00000c9b_sig00001e35 : STD_LOGIC; 
  signal blk00000c9b_sig00001e34 : STD_LOGIC; 
  signal blk00000c9b_sig00001e33 : STD_LOGIC; 
  signal blk00000c9b_sig00001e32 : STD_LOGIC; 
  signal blk00000c9b_sig00001e31 : STD_LOGIC; 
  signal blk00000c9b_sig00001e30 : STD_LOGIC; 
  signal blk00000c9b_sig00001e2f : STD_LOGIC; 
  signal blk00000c9b_sig00001e2e : STD_LOGIC; 
  signal blk00000cb3_sig00001e60 : STD_LOGIC; 
  signal blk00000cb3_sig00001e5f : STD_LOGIC; 
  signal blk00000cb3_sig00001e5e : STD_LOGIC; 
  signal blk00000cb3_sig00001e5d : STD_LOGIC; 
  signal blk00000cb3_sig00001e5c : STD_LOGIC; 
  signal blk00000cb3_sig00001e59 : STD_LOGIC; 
  signal blk00000cb3_sig00001e58 : STD_LOGIC; 
  signal blk00000cb3_sig00001e57 : STD_LOGIC; 
  signal blk00000cb3_sig00001e56 : STD_LOGIC; 
  signal blk00000cb3_sig00001e55 : STD_LOGIC; 
  signal blk00000cb3_sig00001e54 : STD_LOGIC; 
  signal blk00000cb3_sig00001e53 : STD_LOGIC; 
  signal blk00000cb3_sig00001e52 : STD_LOGIC; 
  signal blk00000cb3_sig00001e51 : STD_LOGIC; 
  signal blk00000cb3_sig00001e50 : STD_LOGIC; 
  signal blk00000cb3_sig00001e4f : STD_LOGIC; 
  signal blk00000cb3_sig00001e4e : STD_LOGIC; 
  signal blk00000cb3_sig00001e4d : STD_LOGIC; 
  signal blk00000cb3_sig00001e4c : STD_LOGIC; 
  signal blk00000cb3_sig00001e4b : STD_LOGIC; 
  signal blk00000cb3_sig00001e3f : STD_LOGIC; 
  signal blk00000cb3_sig00001e3e : STD_LOGIC; 
  signal blk00000cb3_sig00001e3d : STD_LOGIC; 
  signal blk00000cd6_blk00000cd7_sig00001e85 : STD_LOGIC; 
  signal blk00000cd6_blk00000cd7_sig00001e84 : STD_LOGIC; 
  signal blk00000cd6_blk00000cd7_sig00001e83 : STD_LOGIC; 
  signal blk00000cd6_blk00000cd7_sig00001e82 : STD_LOGIC; 
  signal blk00000cd6_blk00000cd7_sig00001e81 : STD_LOGIC; 
  signal blk00000cd6_blk00000cd7_sig00001e80 : STD_LOGIC; 
  signal blk00000cd6_blk00000cd7_sig00001e7f : STD_LOGIC; 
  signal blk00000cd6_blk00000cd7_sig00001e7e : STD_LOGIC; 
  signal blk00000ce6_blk00000ce7_sig00001e97 : STD_LOGIC; 
  signal blk00000ce6_blk00000ce7_sig00001e96 : STD_LOGIC; 
  signal blk00000ce6_blk00000ce7_sig00001e95 : STD_LOGIC; 
  signal blk00000cee_sig00001ee5 : STD_LOGIC; 
  signal blk00000cee_sig00001ee4 : STD_LOGIC; 
  signal blk00000cee_sig00001ee3 : STD_LOGIC; 
  signal blk00000cee_sig00001ee2 : STD_LOGIC; 
  signal blk00000cee_sig00001ee1 : STD_LOGIC; 
  signal blk00000cee_sig00001ee0 : STD_LOGIC; 
  signal blk00000cee_sig00001edf : STD_LOGIC; 
  signal blk00000cee_sig00001ede : STD_LOGIC; 
  signal blk00000cee_sig00001edd : STD_LOGIC; 
  signal blk00000cee_sig00001edc : STD_LOGIC; 
  signal blk00000cee_sig00001edb : STD_LOGIC; 
  signal blk00000cee_sig00001eda : STD_LOGIC; 
  signal blk00000cee_sig00001ed9 : STD_LOGIC; 
  signal blk00000cee_sig00001ed8 : STD_LOGIC; 
  signal blk00000cee_sig00001ed7 : STD_LOGIC; 
  signal blk00000cee_sig00001ed6 : STD_LOGIC; 
  signal blk00000cee_sig00001ed5 : STD_LOGIC; 
  signal blk00000cee_sig00001ed4 : STD_LOGIC; 
  signal blk00000cee_sig00001ed3 : STD_LOGIC; 
  signal blk00000cee_sig00001ed2 : STD_LOGIC; 
  signal blk00000cee_sig00001ed1 : STD_LOGIC; 
  signal blk00000cee_sig00001ed0 : STD_LOGIC; 
  signal blk00000cee_sig00001ecf : STD_LOGIC; 
  signal blk00000cee_sig00001ece : STD_LOGIC; 
  signal blk00000cee_sig00001ecd : STD_LOGIC; 
  signal blk00000cee_sig00001ecc : STD_LOGIC; 
  signal blk00000cee_sig00001ecb : STD_LOGIC; 
  signal blk00000cee_sig00001eca : STD_LOGIC; 
  signal blk00000cee_sig00001ec9 : STD_LOGIC; 
  signal blk00000cee_sig00001ec8 : STD_LOGIC; 
  signal blk00000cee_sig00001ec7 : STD_LOGIC; 
  signal blk00000cee_sig00001ec6 : STD_LOGIC; 
  signal blk00000cee_sig00001ec5 : STD_LOGIC; 
  signal blk00000cee_sig00001ec4 : STD_LOGIC; 
  signal blk00000cee_sig00001ec3 : STD_LOGIC; 
  signal blk00000cee_sig00001ec2 : STD_LOGIC; 
  signal blk00000cee_sig00001ec1 : STD_LOGIC; 
  signal blk00000cee_sig00001ec0 : STD_LOGIC; 
  signal blk00000cee_sig00001ebf : STD_LOGIC; 
  signal blk00000d23_sig00001f33 : STD_LOGIC; 
  signal blk00000d23_sig00001f32 : STD_LOGIC; 
  signal blk00000d23_sig00001f31 : STD_LOGIC; 
  signal blk00000d23_sig00001f30 : STD_LOGIC; 
  signal blk00000d23_sig00001f2f : STD_LOGIC; 
  signal blk00000d23_sig00001f2e : STD_LOGIC; 
  signal blk00000d23_sig00001f2d : STD_LOGIC; 
  signal blk00000d23_sig00001f2c : STD_LOGIC; 
  signal blk00000d23_sig00001f2b : STD_LOGIC; 
  signal blk00000d23_sig00001f2a : STD_LOGIC; 
  signal blk00000d23_sig00001f29 : STD_LOGIC; 
  signal blk00000d23_sig00001f28 : STD_LOGIC; 
  signal blk00000d23_sig00001f27 : STD_LOGIC; 
  signal blk00000d23_sig00001f26 : STD_LOGIC; 
  signal blk00000d23_sig00001f25 : STD_LOGIC; 
  signal blk00000d23_sig00001f24 : STD_LOGIC; 
  signal blk00000d23_sig00001f23 : STD_LOGIC; 
  signal blk00000d23_sig00001f22 : STD_LOGIC; 
  signal blk00000d23_sig00001f21 : STD_LOGIC; 
  signal blk00000d23_sig00001f20 : STD_LOGIC; 
  signal blk00000d23_sig00001f1f : STD_LOGIC; 
  signal blk00000d23_sig00001f1e : STD_LOGIC; 
  signal blk00000d23_sig00001f1d : STD_LOGIC; 
  signal blk00000d23_sig00001f1c : STD_LOGIC; 
  signal blk00000d23_sig00001f1b : STD_LOGIC; 
  signal blk00000d23_sig00001f1a : STD_LOGIC; 
  signal blk00000d23_sig00001f19 : STD_LOGIC; 
  signal blk00000d23_sig00001f18 : STD_LOGIC; 
  signal blk00000d23_sig00001f17 : STD_LOGIC; 
  signal blk00000d23_sig00001f16 : STD_LOGIC; 
  signal blk00000d23_sig00001f15 : STD_LOGIC; 
  signal blk00000d23_sig00001f14 : STD_LOGIC; 
  signal blk00000d23_sig00001f13 : STD_LOGIC; 
  signal blk00000d23_sig00001f12 : STD_LOGIC; 
  signal blk00000d23_sig00001f11 : STD_LOGIC; 
  signal blk00000d23_sig00001f10 : STD_LOGIC; 
  signal blk00000d23_sig00001f0f : STD_LOGIC; 
  signal blk00000d23_sig00001f0e : STD_LOGIC; 
  signal blk00000d23_sig00001f0d : STD_LOGIC; 
  signal blk00000d58_blk00000d59_sig00001f44 : STD_LOGIC; 
  signal blk00000d58_blk00000d59_sig00001f43 : STD_LOGIC; 
  signal blk00000d91_blk00000d92_sig00001f86 : STD_LOGIC; 
  signal blk00000d91_blk00000d92_sig00001f85 : STD_LOGIC; 
  signal blk00000d91_blk00000d92_sig00001f84 : STD_LOGIC; 
  signal blk00000d91_blk00000d92_sig00001f83 : STD_LOGIC; 
  signal blk00000d91_blk00000d92_sig00001f82 : STD_LOGIC; 
  signal blk00000d91_blk00000d92_sig00001f81 : STD_LOGIC; 
  signal blk00000d91_blk00000d92_sig00001f80 : STD_LOGIC; 
  signal blk00000d91_blk00000d92_sig00001f7f : STD_LOGIC; 
  signal blk00000d91_blk00000d92_sig00001f7e : STD_LOGIC; 
  signal blk00000d91_blk00000d92_sig00001f7d : STD_LOGIC; 
  signal blk00000d91_blk00000d92_sig00001f7c : STD_LOGIC; 
  signal blk00000d91_blk00000d92_sig00001f7b : STD_LOGIC; 
  signal blk00000d91_blk00000d92_sig00001f7a : STD_LOGIC; 
  signal blk00000dac_blk00000dad_sig00001fc8 : STD_LOGIC; 
  signal blk00000dac_blk00000dad_sig00001fc7 : STD_LOGIC; 
  signal blk00000dac_blk00000dad_sig00001fc6 : STD_LOGIC; 
  signal blk00000dac_blk00000dad_sig00001fc5 : STD_LOGIC; 
  signal blk00000dac_blk00000dad_sig00001fc4 : STD_LOGIC; 
  signal blk00000dac_blk00000dad_sig00001fc3 : STD_LOGIC; 
  signal blk00000dac_blk00000dad_sig00001fc2 : STD_LOGIC; 
  signal blk00000dac_blk00000dad_sig00001fc1 : STD_LOGIC; 
  signal blk00000dac_blk00000dad_sig00001fc0 : STD_LOGIC; 
  signal blk00000dac_blk00000dad_sig00001fbf : STD_LOGIC; 
  signal blk00000dac_blk00000dad_sig00001fbe : STD_LOGIC; 
  signal blk00000dac_blk00000dad_sig00001fbd : STD_LOGIC; 
  signal blk00000dac_blk00000dad_sig00001fbc : STD_LOGIC; 
  signal blk00000dc7_blk00000dc8_sig0000200f : STD_LOGIC; 
  signal blk00000dc7_blk00000dc8_sig0000200e : STD_LOGIC; 
  signal blk00000dc7_blk00000dc8_sig0000200d : STD_LOGIC; 
  signal blk00000dc7_blk00000dc8_sig0000200c : STD_LOGIC; 
  signal blk00000dc7_blk00000dc8_sig0000200b : STD_LOGIC; 
  signal blk00000dc7_blk00000dc8_sig0000200a : STD_LOGIC; 
  signal blk00000dc7_blk00000dc8_sig00002009 : STD_LOGIC; 
  signal blk00000dc7_blk00000dc8_sig00002008 : STD_LOGIC; 
  signal blk00000dc7_blk00000dc8_sig00002007 : STD_LOGIC; 
  signal blk00000dc7_blk00000dc8_sig00002006 : STD_LOGIC; 
  signal blk00000dc7_blk00000dc8_sig00002005 : STD_LOGIC; 
  signal blk00000dc7_blk00000dc8_sig00002004 : STD_LOGIC; 
  signal blk00000dc7_blk00000dc8_sig00002003 : STD_LOGIC; 
  signal blk00000dc7_blk00000dc8_sig00002002 : STD_LOGIC; 
  signal blk00000de4_blk00000de5_sig00002056 : STD_LOGIC; 
  signal blk00000de4_blk00000de5_sig00002055 : STD_LOGIC; 
  signal blk00000de4_blk00000de5_sig00002054 : STD_LOGIC; 
  signal blk00000de4_blk00000de5_sig00002053 : STD_LOGIC; 
  signal blk00000de4_blk00000de5_sig00002052 : STD_LOGIC; 
  signal blk00000de4_blk00000de5_sig00002051 : STD_LOGIC; 
  signal blk00000de4_blk00000de5_sig00002050 : STD_LOGIC; 
  signal blk00000de4_blk00000de5_sig0000204f : STD_LOGIC; 
  signal blk00000de4_blk00000de5_sig0000204e : STD_LOGIC; 
  signal blk00000de4_blk00000de5_sig0000204d : STD_LOGIC; 
  signal blk00000de4_blk00000de5_sig0000204c : STD_LOGIC; 
  signal blk00000de4_blk00000de5_sig0000204b : STD_LOGIC; 
  signal blk00000de4_blk00000de5_sig0000204a : STD_LOGIC; 
  signal blk00000de4_blk00000de5_sig00002049 : STD_LOGIC; 
  signal blk00000e01_blk00000e02_sig00002066 : STD_LOGIC; 
  signal blk00000e01_blk00000e02_sig00002065 : STD_LOGIC; 
  signal blk00000e01_blk00000e02_sig00002064 : STD_LOGIC; 
  signal blk00000e01_blk00000e02_sig00002063 : STD_LOGIC; 
  signal blk00000e09_blk00000e0a_sig00002076 : STD_LOGIC; 
  signal blk00000e09_blk00000e0a_sig00002075 : STD_LOGIC; 
  signal blk00000e09_blk00000e0a_sig00002074 : STD_LOGIC; 
  signal blk00000e09_blk00000e0a_sig00002073 : STD_LOGIC; 
  signal blk00000e11_blk00000e12_sig00002081 : STD_LOGIC; 
  signal blk00000e11_blk00000e12_sig00002080 : STD_LOGIC; 
  signal blk00000e11_blk00000e12_sig0000207f : STD_LOGIC; 
  signal blk00000e17_blk00000e18_sig0000208c : STD_LOGIC; 
  signal blk00000e17_blk00000e18_sig0000208b : STD_LOGIC; 
  signal blk00000e17_blk00000e18_sig0000208a : STD_LOGIC; 
  signal blk00000e1d_blk00000e1e_sig0000209c : STD_LOGIC; 
  signal blk00000e1d_blk00000e1e_sig0000209b : STD_LOGIC; 
  signal blk00000e1d_blk00000e1e_sig0000209a : STD_LOGIC; 
  signal blk00000e1d_blk00000e1e_sig00002099 : STD_LOGIC; 
  signal blk00000e25_blk00000e26_sig000020c0 : STD_LOGIC; 
  signal blk00000e25_blk00000e26_sig000020bf : STD_LOGIC; 
  signal blk00000e25_blk00000e26_sig000020be : STD_LOGIC; 
  signal blk00000e25_blk00000e26_sig000020bd : STD_LOGIC; 
  signal blk00000e25_blk00000e26_sig000020bc : STD_LOGIC; 
  signal blk00000e25_blk00000e26_sig000020bb : STD_LOGIC; 
  signal blk00000e25_blk00000e26_sig000020ba : STD_LOGIC; 
  signal blk00000e25_blk00000e26_sig000020b9 : STD_LOGIC; 
  signal blk00000e35_sig00002116 : STD_LOGIC; 
  signal blk00000e35_sig00002115 : STD_LOGIC; 
  signal blk00000e35_sig00002114 : STD_LOGIC; 
  signal blk00000e35_sig00002113 : STD_LOGIC; 
  signal blk00000e35_sig00002112 : STD_LOGIC; 
  signal blk00000e35_sig00002111 : STD_LOGIC; 
  signal blk00000e35_sig00002110 : STD_LOGIC; 
  signal blk00000e35_sig0000210f : STD_LOGIC; 
  signal blk00000e35_sig0000210e : STD_LOGIC; 
  signal blk00000e35_sig0000210d : STD_LOGIC; 
  signal blk00000e35_sig0000210c : STD_LOGIC; 
  signal blk00000e35_sig0000210b : STD_LOGIC; 
  signal blk00000e35_sig0000210a : STD_LOGIC; 
  signal blk00000e35_sig00002109 : STD_LOGIC; 
  signal blk00000e35_sig00002108 : STD_LOGIC; 
  signal blk00000e35_sig00002107 : STD_LOGIC; 
  signal blk00000e35_sig00002106 : STD_LOGIC; 
  signal blk00000e35_sig00002105 : STD_LOGIC; 
  signal blk00000e35_sig00002104 : STD_LOGIC; 
  signal blk00000e35_sig00002103 : STD_LOGIC; 
  signal blk00000e35_sig00002102 : STD_LOGIC; 
  signal blk00000e35_sig00002101 : STD_LOGIC; 
  signal blk00000e35_sig00002100 : STD_LOGIC; 
  signal blk00000e35_sig000020ff : STD_LOGIC; 
  signal blk00000e35_sig000020fe : STD_LOGIC; 
  signal blk00000e35_sig000020fd : STD_LOGIC; 
  signal blk00000e35_sig000020fc : STD_LOGIC; 
  signal blk00000e35_sig000020fb : STD_LOGIC; 
  signal blk00000e35_sig000020fa : STD_LOGIC; 
  signal blk00000e35_sig000020f9 : STD_LOGIC; 
  signal blk00000e35_sig000020f8 : STD_LOGIC; 
  signal blk00000e35_sig000020f7 : STD_LOGIC; 
  signal blk00000e35_sig000020f6 : STD_LOGIC; 
  signal blk00000e35_sig000020f5 : STD_LOGIC; 
  signal blk00000e35_sig000020f4 : STD_LOGIC; 
  signal blk00000e35_sig000020f3 : STD_LOGIC; 
  signal blk00000e35_sig000020f2 : STD_LOGIC; 
  signal blk00000e35_sig000020f1 : STD_LOGIC; 
  signal blk00000e35_sig000020f0 : STD_LOGIC; 
  signal blk00000e35_sig000020ef : STD_LOGIC; 
  signal blk00000e35_sig000020ee : STD_LOGIC; 
  signal blk00000e35_sig000020ed : STD_LOGIC; 
  signal blk00000e6e_sig0000216c : STD_LOGIC; 
  signal blk00000e6e_sig0000216b : STD_LOGIC; 
  signal blk00000e6e_sig0000216a : STD_LOGIC; 
  signal blk00000e6e_sig00002169 : STD_LOGIC; 
  signal blk00000e6e_sig00002168 : STD_LOGIC; 
  signal blk00000e6e_sig00002167 : STD_LOGIC; 
  signal blk00000e6e_sig00002166 : STD_LOGIC; 
  signal blk00000e6e_sig00002165 : STD_LOGIC; 
  signal blk00000e6e_sig00002164 : STD_LOGIC; 
  signal blk00000e6e_sig00002163 : STD_LOGIC; 
  signal blk00000e6e_sig00002162 : STD_LOGIC; 
  signal blk00000e6e_sig00002161 : STD_LOGIC; 
  signal blk00000e6e_sig00002160 : STD_LOGIC; 
  signal blk00000e6e_sig0000215f : STD_LOGIC; 
  signal blk00000e6e_sig0000215e : STD_LOGIC; 
  signal blk00000e6e_sig0000215d : STD_LOGIC; 
  signal blk00000e6e_sig0000215c : STD_LOGIC; 
  signal blk00000e6e_sig0000215b : STD_LOGIC; 
  signal blk00000e6e_sig0000215a : STD_LOGIC; 
  signal blk00000e6e_sig00002159 : STD_LOGIC; 
  signal blk00000e6e_sig00002158 : STD_LOGIC; 
  signal blk00000e6e_sig00002157 : STD_LOGIC; 
  signal blk00000e6e_sig00002156 : STD_LOGIC; 
  signal blk00000e6e_sig00002155 : STD_LOGIC; 
  signal blk00000e6e_sig00002154 : STD_LOGIC; 
  signal blk00000e6e_sig00002153 : STD_LOGIC; 
  signal blk00000e6e_sig00002152 : STD_LOGIC; 
  signal blk00000e6e_sig00002151 : STD_LOGIC; 
  signal blk00000e6e_sig00002150 : STD_LOGIC; 
  signal blk00000e6e_sig0000214f : STD_LOGIC; 
  signal blk00000e6e_sig0000214e : STD_LOGIC; 
  signal blk00000e6e_sig0000214d : STD_LOGIC; 
  signal blk00000e6e_sig0000214c : STD_LOGIC; 
  signal blk00000e6e_sig0000214b : STD_LOGIC; 
  signal blk00000e6e_sig0000214a : STD_LOGIC; 
  signal blk00000e6e_sig00002149 : STD_LOGIC; 
  signal blk00000e6e_sig00002148 : STD_LOGIC; 
  signal blk00000e6e_sig00002147 : STD_LOGIC; 
  signal blk00000e6e_sig00002146 : STD_LOGIC; 
  signal blk00000e6e_sig00002145 : STD_LOGIC; 
  signal blk00000e6e_sig00002144 : STD_LOGIC; 
  signal blk00000e6e_sig00002143 : STD_LOGIC; 
  signal blk00000ea7_blk00000ea8_sig0000217d : STD_LOGIC; 
  signal blk00000ea7_blk00000ea8_sig0000217c : STD_LOGIC; 
  signal blk00000eac_blk00000ead_sig0000218e : STD_LOGIC; 
  signal blk00000eac_blk00000ead_sig0000218d : STD_LOGIC; 
  signal blk00000fbf_sig000021cf : STD_LOGIC; 
  signal blk00000fc2_blk00000fc3_sig000021f4 : STD_LOGIC; 
  signal blk00000fc2_blk00000fc3_sig000021f3 : STD_LOGIC; 
  signal blk00000fc2_blk00000fc3_sig000021f2 : STD_LOGIC; 
  signal blk00000fc2_blk00000fc3_sig000021f1 : STD_LOGIC; 
  signal blk00000fc2_blk00000fc3_sig000021f0 : STD_LOGIC; 
  signal blk00000fc2_blk00000fc3_sig000021ef : STD_LOGIC; 
  signal blk00000fc2_blk00000fc3_sig000021ee : STD_LOGIC; 
  signal blk00000fc2_blk00000fc3_sig000021ed : STD_LOGIC; 
  signal blk00000fd8_blk00000fd9_sig00002205 : STD_LOGIC; 
  signal blk00000fd8_blk00000fd9_sig00002204 : STD_LOGIC; 
  signal NLW_blk0000040d_O_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk0000042a_O_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000655_PATTERNBDETECT_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000655_PATTERNDETECT_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000655_OVERFLOW_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000655_UNDERFLOW_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000655_CARRYCASCOUT_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000655_MULTSIGNOUT_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000655_PCOUT_47_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000655_PCOUT_46_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000655_PCOUT_45_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000655_PCOUT_44_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000655_PCOUT_43_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000655_PCOUT_42_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000655_PCOUT_41_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000655_PCOUT_40_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000655_PCOUT_39_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000655_PCOUT_38_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000655_PCOUT_37_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000655_PCOUT_36_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000655_PCOUT_35_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000655_PCOUT_34_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000655_PCOUT_33_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000655_PCOUT_32_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000655_PCOUT_31_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000655_PCOUT_30_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000655_PCOUT_29_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000655_PCOUT_28_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000655_PCOUT_27_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000655_PCOUT_26_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000655_PCOUT_25_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000655_PCOUT_24_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000655_PCOUT_23_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000655_PCOUT_22_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000655_PCOUT_21_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000655_PCOUT_20_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000655_PCOUT_19_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000655_PCOUT_18_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000655_PCOUT_17_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000655_PCOUT_16_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000655_PCOUT_15_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000655_PCOUT_14_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000655_PCOUT_13_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000655_PCOUT_12_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000655_PCOUT_11_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000655_PCOUT_10_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000655_PCOUT_9_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000655_PCOUT_8_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000655_PCOUT_7_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000655_PCOUT_6_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000655_PCOUT_5_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000655_PCOUT_4_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000655_PCOUT_3_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000655_PCOUT_2_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000655_PCOUT_1_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000655_PCOUT_0_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000655_P_47_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000655_P_46_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000655_P_45_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000655_P_44_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000655_P_43_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000655_BCOUT_17_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000655_BCOUT_16_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000655_BCOUT_15_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000655_BCOUT_14_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000655_BCOUT_13_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000655_BCOUT_12_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000655_BCOUT_11_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000655_BCOUT_10_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000655_BCOUT_9_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000655_BCOUT_8_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000655_BCOUT_7_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000655_BCOUT_6_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000655_BCOUT_5_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000655_BCOUT_4_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000655_BCOUT_3_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000655_BCOUT_2_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000655_BCOUT_1_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000655_BCOUT_0_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000655_ACOUT_29_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000655_ACOUT_28_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000655_ACOUT_27_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000655_ACOUT_26_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000655_ACOUT_25_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000655_ACOUT_24_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000655_ACOUT_23_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000655_ACOUT_22_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000655_ACOUT_21_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000655_ACOUT_20_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000655_ACOUT_19_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000655_ACOUT_18_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000655_ACOUT_17_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000655_ACOUT_16_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000655_ACOUT_15_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000655_ACOUT_14_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000655_ACOUT_13_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000655_ACOUT_12_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000655_ACOUT_11_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000655_ACOUT_10_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000655_ACOUT_9_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000655_ACOUT_8_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000655_ACOUT_7_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000655_ACOUT_6_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000655_ACOUT_5_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000655_ACOUT_4_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000655_ACOUT_3_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000655_ACOUT_2_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000655_ACOUT_1_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000655_ACOUT_0_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000655_CARRYOUT_3_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000655_CARRYOUT_2_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000655_CARRYOUT_1_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000655_CARRYOUT_0_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000656_PATTERNBDETECT_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000656_PATTERNDETECT_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000656_OVERFLOW_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000656_UNDERFLOW_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000656_CARRYCASCOUT_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000656_MULTSIGNOUT_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000656_PCOUT_47_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000656_PCOUT_46_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000656_PCOUT_45_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000656_PCOUT_44_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000656_PCOUT_43_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000656_PCOUT_42_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000656_PCOUT_41_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000656_PCOUT_40_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000656_PCOUT_39_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000656_PCOUT_38_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000656_PCOUT_37_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000656_PCOUT_36_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000656_PCOUT_35_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000656_PCOUT_34_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000656_PCOUT_33_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000656_PCOUT_32_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000656_PCOUT_31_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000656_PCOUT_30_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000656_PCOUT_29_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000656_PCOUT_28_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000656_PCOUT_27_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000656_PCOUT_26_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000656_PCOUT_25_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000656_PCOUT_24_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000656_PCOUT_23_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000656_PCOUT_22_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000656_PCOUT_21_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000656_PCOUT_20_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000656_PCOUT_19_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000656_PCOUT_18_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000656_PCOUT_17_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000656_PCOUT_16_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000656_PCOUT_15_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000656_PCOUT_14_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000656_PCOUT_13_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000656_PCOUT_12_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000656_PCOUT_11_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000656_PCOUT_10_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000656_PCOUT_9_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000656_PCOUT_8_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000656_PCOUT_7_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000656_PCOUT_6_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000656_PCOUT_5_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000656_PCOUT_4_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000656_PCOUT_3_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000656_PCOUT_2_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000656_PCOUT_1_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000656_PCOUT_0_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000656_P_47_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000656_P_46_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000656_P_45_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000656_P_44_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000656_P_43_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000656_BCOUT_17_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000656_BCOUT_16_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000656_BCOUT_15_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000656_BCOUT_14_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000656_BCOUT_13_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000656_BCOUT_12_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000656_BCOUT_11_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000656_BCOUT_10_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000656_BCOUT_9_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000656_BCOUT_8_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000656_BCOUT_7_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000656_BCOUT_6_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000656_BCOUT_5_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000656_BCOUT_4_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000656_BCOUT_3_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000656_BCOUT_2_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000656_BCOUT_1_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000656_BCOUT_0_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000656_ACOUT_29_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000656_ACOUT_28_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000656_ACOUT_27_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000656_ACOUT_26_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000656_ACOUT_25_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000656_ACOUT_24_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000656_ACOUT_23_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000656_ACOUT_22_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000656_ACOUT_21_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000656_ACOUT_20_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000656_ACOUT_19_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000656_ACOUT_18_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000656_ACOUT_17_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000656_ACOUT_16_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000656_ACOUT_15_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000656_ACOUT_14_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000656_ACOUT_13_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000656_ACOUT_12_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000656_ACOUT_11_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000656_ACOUT_10_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000656_ACOUT_9_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000656_ACOUT_8_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000656_ACOUT_7_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000656_ACOUT_6_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000656_ACOUT_5_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000656_ACOUT_4_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000656_ACOUT_3_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000656_ACOUT_2_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000656_ACOUT_1_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000656_ACOUT_0_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000656_CARRYOUT_3_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000656_CARRYOUT_2_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000656_CARRYOUT_1_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000656_CARRYOUT_0_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000657_PATTERNBDETECT_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000657_PATTERNDETECT_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000657_OVERFLOW_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000657_UNDERFLOW_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000657_CARRYCASCOUT_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000657_MULTSIGNOUT_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000657_PCOUT_47_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000657_PCOUT_46_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000657_PCOUT_45_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000657_PCOUT_44_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000657_PCOUT_43_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000657_PCOUT_42_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000657_PCOUT_41_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000657_PCOUT_40_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000657_PCOUT_39_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000657_PCOUT_38_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000657_PCOUT_37_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000657_PCOUT_36_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000657_PCOUT_35_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000657_PCOUT_34_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000657_PCOUT_33_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000657_PCOUT_32_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000657_PCOUT_31_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000657_PCOUT_30_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000657_PCOUT_29_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000657_PCOUT_28_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000657_PCOUT_27_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000657_PCOUT_26_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000657_PCOUT_25_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000657_PCOUT_24_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000657_PCOUT_23_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000657_PCOUT_22_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000657_PCOUT_21_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000657_PCOUT_20_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000657_PCOUT_19_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000657_PCOUT_18_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000657_PCOUT_17_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000657_PCOUT_16_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000657_PCOUT_15_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000657_PCOUT_14_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000657_PCOUT_13_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000657_PCOUT_12_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000657_PCOUT_11_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000657_PCOUT_10_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000657_PCOUT_9_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000657_PCOUT_8_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000657_PCOUT_7_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000657_PCOUT_6_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000657_PCOUT_5_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000657_PCOUT_4_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000657_PCOUT_3_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000657_PCOUT_2_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000657_PCOUT_1_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000657_PCOUT_0_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000657_P_47_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000657_P_46_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000657_P_45_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000657_P_44_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000657_P_43_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000657_BCOUT_17_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000657_BCOUT_16_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000657_BCOUT_15_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000657_BCOUT_14_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000657_BCOUT_13_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000657_BCOUT_12_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000657_BCOUT_11_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000657_BCOUT_10_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000657_BCOUT_9_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000657_BCOUT_8_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000657_BCOUT_7_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000657_BCOUT_6_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000657_BCOUT_5_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000657_BCOUT_4_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000657_BCOUT_3_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000657_BCOUT_2_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000657_BCOUT_1_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000657_BCOUT_0_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000657_ACOUT_29_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000657_ACOUT_28_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000657_ACOUT_27_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000657_ACOUT_26_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000657_ACOUT_25_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000657_ACOUT_24_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000657_ACOUT_23_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000657_ACOUT_22_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000657_ACOUT_21_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000657_ACOUT_20_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000657_ACOUT_19_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000657_ACOUT_18_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000657_ACOUT_17_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000657_ACOUT_16_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000657_ACOUT_15_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000657_ACOUT_14_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000657_ACOUT_13_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000657_ACOUT_12_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000657_ACOUT_11_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000657_ACOUT_10_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000657_ACOUT_9_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000657_ACOUT_8_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000657_ACOUT_7_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000657_ACOUT_6_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000657_ACOUT_5_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000657_ACOUT_4_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000657_ACOUT_3_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000657_ACOUT_2_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000657_ACOUT_1_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000657_ACOUT_0_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000657_CARRYOUT_3_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000657_CARRYOUT_2_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000657_CARRYOUT_1_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000657_CARRYOUT_0_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk0000077e_Q_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk0000077f_Q_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000780_Q_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000781_Q_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000782_Q_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000783_Q_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000784_Q_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000785_Q_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000792_Q_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000793_Q_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000794_Q_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk000007ac_Q_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk000007ad_Q_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk000007ae_Q_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk000007af_Q_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk000007b0_Q_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk000007b1_Q_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk000007b2_Q_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk000007b3_Q_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk000007c0_Q_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk000007c1_Q_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk000007c2_Q_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk000007c3_Q_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk000007c4_Q_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk000007c5_Q_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk000007d2_Q_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk000007d3_Q_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk000007d4_Q_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk000007d5_Q_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk000007d6_Q_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk000007d7_Q_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk000007d8_Q_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk000007d9_Q_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk000007f1_Q_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk000007f2_Q_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk000007f3_Q_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000800_Q_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000801_Q_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000802_Q_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000803_Q_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000804_Q_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000805_Q_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000806_Q_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000807_Q_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000917_PATTERNBDETECT_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000917_PATTERNDETECT_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000917_OVERFLOW_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000917_UNDERFLOW_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000917_CARRYCASCOUT_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000917_MULTSIGNOUT_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000917_PCOUT_47_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000917_PCOUT_46_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000917_PCOUT_45_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000917_PCOUT_44_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000917_PCOUT_43_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000917_PCOUT_42_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000917_PCOUT_41_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000917_PCOUT_40_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000917_PCOUT_39_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000917_PCOUT_38_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000917_PCOUT_37_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000917_PCOUT_36_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000917_PCOUT_35_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000917_PCOUT_34_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000917_PCOUT_33_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000917_PCOUT_32_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000917_PCOUT_31_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000917_PCOUT_30_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000917_PCOUT_29_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000917_PCOUT_28_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000917_PCOUT_27_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000917_PCOUT_26_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000917_PCOUT_25_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000917_PCOUT_24_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000917_PCOUT_23_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000917_PCOUT_22_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000917_PCOUT_21_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000917_PCOUT_20_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000917_PCOUT_19_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000917_PCOUT_18_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000917_PCOUT_17_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000917_PCOUT_16_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000917_PCOUT_15_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000917_PCOUT_14_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000917_PCOUT_13_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000917_PCOUT_12_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000917_PCOUT_11_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000917_PCOUT_10_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000917_PCOUT_9_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000917_PCOUT_8_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000917_PCOUT_7_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000917_PCOUT_6_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000917_PCOUT_5_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000917_PCOUT_4_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000917_PCOUT_3_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000917_PCOUT_2_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000917_PCOUT_1_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000917_PCOUT_0_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000917_P_47_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000917_P_46_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000917_P_45_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000917_P_44_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000917_P_43_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000917_BCOUT_17_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000917_BCOUT_16_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000917_BCOUT_15_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000917_BCOUT_14_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000917_BCOUT_13_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000917_BCOUT_12_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000917_BCOUT_11_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000917_BCOUT_10_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000917_BCOUT_9_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000917_BCOUT_8_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000917_BCOUT_7_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000917_BCOUT_6_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000917_BCOUT_5_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000917_BCOUT_4_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000917_BCOUT_3_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000917_BCOUT_2_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000917_BCOUT_1_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000917_BCOUT_0_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000917_ACOUT_29_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000917_ACOUT_28_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000917_ACOUT_27_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000917_ACOUT_26_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000917_ACOUT_25_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000917_ACOUT_24_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000917_ACOUT_23_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000917_ACOUT_22_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000917_ACOUT_21_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000917_ACOUT_20_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000917_ACOUT_19_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000917_ACOUT_18_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000917_ACOUT_17_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000917_ACOUT_16_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000917_ACOUT_15_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000917_ACOUT_14_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000917_ACOUT_13_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000917_ACOUT_12_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000917_ACOUT_11_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000917_ACOUT_10_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000917_ACOUT_9_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000917_ACOUT_8_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000917_ACOUT_7_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000917_ACOUT_6_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000917_ACOUT_5_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000917_ACOUT_4_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000917_ACOUT_3_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000917_ACOUT_2_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000917_ACOUT_1_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000917_ACOUT_0_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000917_CARRYOUT_3_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000917_CARRYOUT_2_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000917_CARRYOUT_1_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000917_CARRYOUT_0_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000918_PATTERNBDETECT_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000918_PATTERNDETECT_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000918_OVERFLOW_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000918_UNDERFLOW_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000918_CARRYCASCOUT_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000918_MULTSIGNOUT_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000918_PCOUT_47_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000918_PCOUT_46_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000918_PCOUT_45_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000918_PCOUT_44_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000918_PCOUT_43_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000918_PCOUT_42_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000918_PCOUT_41_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000918_PCOUT_40_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000918_PCOUT_39_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000918_PCOUT_38_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000918_PCOUT_37_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000918_PCOUT_36_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000918_PCOUT_35_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000918_PCOUT_34_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000918_PCOUT_33_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000918_PCOUT_32_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000918_PCOUT_31_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000918_PCOUT_30_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000918_PCOUT_29_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000918_PCOUT_28_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000918_PCOUT_27_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000918_PCOUT_26_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000918_PCOUT_25_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000918_PCOUT_24_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000918_PCOUT_23_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000918_PCOUT_22_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000918_PCOUT_21_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000918_PCOUT_20_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000918_PCOUT_19_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000918_PCOUT_18_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000918_PCOUT_17_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000918_PCOUT_16_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000918_PCOUT_15_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000918_PCOUT_14_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000918_PCOUT_13_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000918_PCOUT_12_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000918_PCOUT_11_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000918_PCOUT_10_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000918_PCOUT_9_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000918_PCOUT_8_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000918_PCOUT_7_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000918_PCOUT_6_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000918_PCOUT_5_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000918_PCOUT_4_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000918_PCOUT_3_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000918_PCOUT_2_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000918_PCOUT_1_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000918_PCOUT_0_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000918_P_47_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000918_P_46_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000918_P_45_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000918_P_44_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000918_P_43_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000918_BCOUT_17_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000918_BCOUT_16_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000918_BCOUT_15_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000918_BCOUT_14_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000918_BCOUT_13_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000918_BCOUT_12_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000918_BCOUT_11_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000918_BCOUT_10_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000918_BCOUT_9_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000918_BCOUT_8_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000918_BCOUT_7_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000918_BCOUT_6_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000918_BCOUT_5_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000918_BCOUT_4_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000918_BCOUT_3_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000918_BCOUT_2_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000918_BCOUT_1_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000918_BCOUT_0_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000918_ACOUT_29_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000918_ACOUT_28_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000918_ACOUT_27_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000918_ACOUT_26_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000918_ACOUT_25_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000918_ACOUT_24_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000918_ACOUT_23_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000918_ACOUT_22_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000918_ACOUT_21_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000918_ACOUT_20_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000918_ACOUT_19_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000918_ACOUT_18_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000918_ACOUT_17_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000918_ACOUT_16_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000918_ACOUT_15_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000918_ACOUT_14_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000918_ACOUT_13_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000918_ACOUT_12_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000918_ACOUT_11_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000918_ACOUT_10_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000918_ACOUT_9_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000918_ACOUT_8_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000918_ACOUT_7_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000918_ACOUT_6_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000918_ACOUT_5_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000918_ACOUT_4_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000918_ACOUT_3_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000918_ACOUT_2_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000918_ACOUT_1_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000918_ACOUT_0_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000918_CARRYOUT_3_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000918_CARRYOUT_2_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000918_CARRYOUT_1_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000918_CARRYOUT_0_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000919_PATTERNBDETECT_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000919_PATTERNDETECT_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000919_OVERFLOW_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000919_UNDERFLOW_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000919_CARRYCASCOUT_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000919_MULTSIGNOUT_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000919_PCOUT_47_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000919_PCOUT_46_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000919_PCOUT_45_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000919_PCOUT_44_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000919_PCOUT_43_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000919_PCOUT_42_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000919_PCOUT_41_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000919_PCOUT_40_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000919_PCOUT_39_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000919_PCOUT_38_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000919_PCOUT_37_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000919_PCOUT_36_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000919_PCOUT_35_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000919_PCOUT_34_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000919_PCOUT_33_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000919_PCOUT_32_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000919_PCOUT_31_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000919_PCOUT_30_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000919_PCOUT_29_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000919_PCOUT_28_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000919_PCOUT_27_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000919_PCOUT_26_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000919_PCOUT_25_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000919_PCOUT_24_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000919_PCOUT_23_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000919_PCOUT_22_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000919_PCOUT_21_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000919_PCOUT_20_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000919_PCOUT_19_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000919_PCOUT_18_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000919_PCOUT_17_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000919_PCOUT_16_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000919_PCOUT_15_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000919_PCOUT_14_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000919_PCOUT_13_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000919_PCOUT_12_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000919_PCOUT_11_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000919_PCOUT_10_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000919_PCOUT_9_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000919_PCOUT_8_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000919_PCOUT_7_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000919_PCOUT_6_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000919_PCOUT_5_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000919_PCOUT_4_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000919_PCOUT_3_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000919_PCOUT_2_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000919_PCOUT_1_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000919_PCOUT_0_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000919_P_47_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000919_P_46_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000919_P_45_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000919_P_44_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000919_P_43_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000919_BCOUT_17_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000919_BCOUT_16_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000919_BCOUT_15_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000919_BCOUT_14_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000919_BCOUT_13_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000919_BCOUT_12_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000919_BCOUT_11_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000919_BCOUT_10_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000919_BCOUT_9_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000919_BCOUT_8_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000919_BCOUT_7_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000919_BCOUT_6_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000919_BCOUT_5_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000919_BCOUT_4_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000919_BCOUT_3_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000919_BCOUT_2_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000919_BCOUT_1_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000919_BCOUT_0_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000919_ACOUT_29_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000919_ACOUT_28_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000919_ACOUT_27_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000919_ACOUT_26_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000919_ACOUT_25_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000919_ACOUT_24_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000919_ACOUT_23_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000919_ACOUT_22_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000919_ACOUT_21_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000919_ACOUT_20_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000919_ACOUT_19_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000919_ACOUT_18_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000919_ACOUT_17_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000919_ACOUT_16_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000919_ACOUT_15_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000919_ACOUT_14_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000919_ACOUT_13_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000919_ACOUT_12_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000919_ACOUT_11_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000919_ACOUT_10_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000919_ACOUT_9_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000919_ACOUT_8_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000919_ACOUT_7_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000919_ACOUT_6_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000919_ACOUT_5_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000919_ACOUT_4_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000919_ACOUT_3_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000919_ACOUT_2_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000919_ACOUT_1_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000919_ACOUT_0_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000919_CARRYOUT_3_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000919_CARRYOUT_2_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000919_CARRYOUT_1_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000919_CARRYOUT_0_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000b73_O_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000b90_O_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000ecb_O_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000ee8_O_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000f8c_Q_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000f8d_Q_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000f8e_Q_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000f9b_Q_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000f9c_Q_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000fae_Q_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000faf_Q_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000fb0_Q_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000fbd_Q_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000fbe_Q_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00001256_Q15_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00001258_Q15_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk0000125a_Q15_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk0000125c_Q15_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk0000125e_Q15_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00001260_Q15_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00001262_Q15_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00001264_Q15_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00001266_Q15_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00001268_Q15_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk0000126a_Q15_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk0000126c_Q15_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk0000126e_Q15_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00001270_Q15_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00001272_Q15_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00001274_Q15_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00001276_Q15_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00001278_Q15_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk0000127a_Q15_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk0000127c_Q15_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk0000127e_Q15_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00001280_Q15_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00001282_Q15_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00001284_Q15_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00001286_Q15_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00001288_Q15_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk0000128a_Q15_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk0000128c_Q15_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk0000128e_Q15_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00001290_Q15_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00001292_Q15_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00001294_Q15_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00001296_Q15_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00001298_Q15_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk0000129a_Q15_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk0000129c_Q15_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk0000129e_Q15_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk000012a0_Q15_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk000012a2_Q15_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk000012a4_Q15_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk000012a6_Q15_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk000012a8_Q15_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk000012aa_Q15_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk000012ac_Q15_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk000012ae_Q15_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk000012b0_Q15_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk000012b2_Q15_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk000012b4_Q15_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk000012b6_Q15_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk000012b8_Q15_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk000012ba_Q15_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk000012bc_Q15_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk000012be_Q15_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk000012c0_Q15_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk000012c2_Q15_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk000012c4_Q15_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk000012c6_Q15_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk000012c8_Q15_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk000012ca_Q15_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk000012cc_Q15_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk000012ce_Q15_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk000012d0_Q15_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk000012d2_Q15_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk000012d4_Q15_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk000012d6_Q15_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk000012d8_Q15_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk000012da_Q15_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk000012dc_Q15_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk000012de_Q15_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk000012e0_Q15_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk000012e2_Q15_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk000012e4_Q15_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk000012e6_Q15_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk000012e8_Q15_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk000012ea_Q15_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk000012ec_Q15_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk000012ee_Q15_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk000012f0_Q15_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk000012f2_Q15_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk000012f4_Q15_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk000012f6_Q15_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk000012f8_Q15_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk000012fa_Q15_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk000012fc_Q15_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk000012fe_Q15_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00001300_Q15_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00001302_Q15_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00001304_Q15_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00001306_Q15_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00001308_Q15_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk0000130a_Q15_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk0000130c_Q15_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk0000130e_Q15_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00001310_Q15_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00001312_Q15_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00001314_Q15_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00001316_Q15_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00001318_Q15_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk0000131a_Q15_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk0000131c_Q15_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk0000131e_Q15_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00001320_Q15_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00001322_Q15_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00001324_Q15_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00001326_Q15_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00001328_Q15_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk0000132a_Q15_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk0000132c_Q15_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk0000132e_Q15_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00001330_Q15_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00001332_Q15_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00001334_Q15_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00001336_Q15_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00001338_Q15_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk0000133a_Q15_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk0000133c_Q15_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk0000133e_Q15_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00001340_Q15_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00001342_Q15_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00001344_Q15_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00001346_Q15_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00001348_Q15_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk0000134a_Q15_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk0000134c_Q15_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk0000134e_Q15_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00001350_Q15_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00001352_Q15_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00001354_Q15_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00001356_Q15_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00001358_Q15_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000065_blk00000066_blk0000007f_Q15_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000065_blk00000066_blk0000007d_Q15_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000065_blk00000066_blk0000007b_Q15_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000065_blk00000066_blk00000079_Q15_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000065_blk00000066_blk00000077_Q15_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000065_blk00000066_blk00000075_Q15_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000065_blk00000066_blk00000073_Q15_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000065_blk00000066_blk00000071_Q15_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000065_blk00000066_blk0000006f_Q15_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000065_blk00000066_blk0000006d_Q15_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000065_blk00000066_blk0000006b_Q15_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000065_blk00000066_blk00000069_Q15_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000081_blk00000082_blk0000009b_Q15_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000081_blk00000082_blk00000099_Q15_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000081_blk00000082_blk00000097_Q15_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000081_blk00000082_blk00000095_Q15_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000081_blk00000082_blk00000093_Q15_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000081_blk00000082_blk00000091_Q15_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000081_blk00000082_blk0000008f_Q15_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000081_blk00000082_blk0000008d_Q15_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000081_blk00000082_blk0000008b_Q15_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000081_blk00000082_blk00000089_Q15_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000081_blk00000082_blk00000087_Q15_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000081_blk00000082_blk00000085_Q15_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk0000017b_blk0000017c_blk0000017f_Q15_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000181_blk00000182_blk00000185_Q15_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000187_blk00000188_blk0000018b_Q15_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk0000018d_blk0000018e_blk00000191_Q15_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000193_blk00000194_blk00000199_Q15_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000193_blk00000194_blk00000197_Q15_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk000001fa_blk000001fb_blk000001fe_Q15_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000200_blk00000201_blk0000021a_Q15_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000200_blk00000201_blk00000218_Q15_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000200_blk00000201_blk00000216_Q15_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000200_blk00000201_blk00000214_Q15_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000200_blk00000201_blk00000212_Q15_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000200_blk00000201_blk00000210_Q15_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000200_blk00000201_blk0000020e_Q15_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000200_blk00000201_blk0000020c_Q15_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000200_blk00000201_blk0000020a_Q15_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000200_blk00000201_blk00000208_Q15_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000200_blk00000201_blk00000206_Q15_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000200_blk00000201_blk00000204_Q15_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk0000021c_blk0000021d_blk00000236_Q15_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk0000021c_blk0000021d_blk00000234_Q15_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk0000021c_blk0000021d_blk00000232_Q15_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk0000021c_blk0000021d_blk00000230_Q15_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk0000021c_blk0000021d_blk0000022e_Q15_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk0000021c_blk0000021d_blk0000022c_Q15_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk0000021c_blk0000021d_blk0000022a_Q15_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk0000021c_blk0000021d_blk00000228_Q15_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk0000021c_blk0000021d_blk00000226_Q15_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk0000021c_blk0000021d_blk00000224_Q15_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk0000021c_blk0000021d_blk00000222_Q15_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk0000021c_blk0000021d_blk00000220_Q15_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000287_blk00000288_blk000002bd_Q31_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000287_blk00000288_blk000002bb_Q31_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000287_blk00000288_blk000002b9_Q31_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000287_blk00000288_blk000002b7_Q31_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000287_blk00000288_blk000002b5_Q31_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000287_blk00000288_blk000002b3_Q31_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000287_blk00000288_blk000002b1_Q31_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000287_blk00000288_blk000002af_Q31_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000287_blk00000288_blk000002ad_Q31_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000287_blk00000288_blk000002ab_Q31_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000287_blk00000288_blk000002a9_Q31_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000287_blk00000288_blk000002a7_Q31_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000287_blk00000288_blk000002a5_Q31_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000287_blk00000288_blk000002a3_Q31_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000287_blk00000288_blk000002a1_Q31_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000287_blk00000288_blk0000029f_Q31_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000287_blk00000288_blk0000029d_Q31_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000287_blk00000288_blk0000029b_Q31_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000287_blk00000288_blk00000299_Q31_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000287_blk00000288_blk00000297_Q31_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000287_blk00000288_blk00000295_Q31_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000287_blk00000288_blk00000293_Q31_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000287_blk00000288_blk00000291_Q31_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000287_blk00000288_blk0000028f_Q31_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000287_blk00000288_blk0000028d_Q31_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000287_blk00000288_blk0000028b_Q31_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk000003bb_blk000003bc_blk000003be_Q31_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk000003c0_blk000003c1_blk000003cd_Q31_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk000003c0_blk000003c1_blk000003cb_Q31_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk000003c0_blk000003c1_blk000003c9_Q31_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk000003c0_blk000003c1_blk000003c7_Q31_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk000003c0_blk000003c1_blk000003c5_Q31_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk000003c0_blk000003c1_blk000003c3_Q31_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk000003cf_blk000003d0_blk000003d3_Q31_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk000003d5_blk000003d6_blk000003d9_Q15_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk000003db_blk000003dc_blk000003de_Q31_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk000003e0_blk000003e1_blk000003e6_Q31_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk000003e0_blk000003e1_blk000003e4_Q31_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk000003e8_blk000003e9_blk000003f1_Q31_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk000003e8_blk000003e9_blk000003ef_Q31_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk000003e8_blk000003e9_blk000003ed_Q31_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk000003e8_blk000003e9_blk000003eb_Q31_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk000004a0_blk000004a1_blk000004a3_Q15_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk000004a5_blk000004a6_blk000004a8_Q15_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk000004aa_blk000004ab_blk000004ad_Q15_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk000004af_blk000004b0_blk000004b2_Q15_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk000004b4_blk000004b5_blk000004b8_Q15_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk000004ba_blk000004bb_blk000004d8_Q15_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk000004ba_blk000004bb_blk000004d6_Q15_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk000004ba_blk000004bb_blk000004d4_Q15_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk000004ba_blk000004bb_blk000004d2_Q15_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk000004ba_blk000004bb_blk000004d0_Q15_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk000004ba_blk000004bb_blk000004ce_Q15_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk000004ba_blk000004bb_blk000004cc_Q15_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk000004ba_blk000004bb_blk000004ca_Q15_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk000004ba_blk000004bb_blk000004c8_Q15_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk000004ba_blk000004bb_blk000004c6_Q15_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk000004ba_blk000004bb_blk000004c4_Q15_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk000004ba_blk000004bb_blk000004c2_Q15_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk000004ba_blk000004bb_blk000004c0_Q15_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk000004ba_blk000004bb_blk000004be_Q15_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk000004da_blk000004db_blk000004f8_Q15_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk000004da_blk000004db_blk000004f6_Q15_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk000004da_blk000004db_blk000004f4_Q15_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk000004da_blk000004db_blk000004f2_Q15_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk000004da_blk000004db_blk000004f0_Q15_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk000004da_blk000004db_blk000004ee_Q15_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk000004da_blk000004db_blk000004ec_Q15_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk000004da_blk000004db_blk000004ea_Q15_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk000004da_blk000004db_blk000004e8_Q15_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk000004da_blk000004db_blk000004e6_Q15_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk000004da_blk000004db_blk000004e4_Q15_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk000004da_blk000004db_blk000004e2_Q15_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk000004da_blk000004db_blk000004e0_Q15_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk000004da_blk000004db_blk000004de_Q15_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk000004fa_blk000004fb_blk00000518_Q15_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk000004fa_blk000004fb_blk00000516_Q15_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk000004fa_blk000004fb_blk00000514_Q15_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk000004fa_blk000004fb_blk00000512_Q15_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk000004fa_blk000004fb_blk00000510_Q15_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk000004fa_blk000004fb_blk0000050e_Q15_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk000004fa_blk000004fb_blk0000050c_Q15_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk000004fa_blk000004fb_blk0000050a_Q15_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk000004fa_blk000004fb_blk00000508_Q15_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk000004fa_blk000004fb_blk00000506_Q15_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk000004fa_blk000004fb_blk00000504_Q15_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk000004fa_blk000004fb_blk00000502_Q15_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk000004fa_blk000004fb_blk00000500_Q15_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk000004fa_blk000004fb_blk000004fe_Q15_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk0000051a_blk0000051b_blk00000538_Q15_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk0000051a_blk0000051b_blk00000536_Q15_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk0000051a_blk0000051b_blk00000534_Q15_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk0000051a_blk0000051b_blk00000532_Q15_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk0000051a_blk0000051b_blk00000530_Q15_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk0000051a_blk0000051b_blk0000052e_Q15_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk0000051a_blk0000051b_blk0000052c_Q15_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk0000051a_blk0000051b_blk0000052a_Q15_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk0000051a_blk0000051b_blk00000528_Q15_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk0000051a_blk0000051b_blk00000526_Q15_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk0000051a_blk0000051b_blk00000524_Q15_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk0000051a_blk0000051b_blk00000522_Q15_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk0000051a_blk0000051b_blk00000520_Q15_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk0000051a_blk0000051b_blk0000051e_Q15_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk000005ac_blk000005ad_blk000005ba_Q31_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk000005ac_blk000005ad_blk000005b8_Q31_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk000005ac_blk000005ad_blk000005b6_Q31_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk000005ac_blk000005ad_blk000005b4_Q31_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk000005ac_blk000005ad_blk000005b2_Q31_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk000005ac_blk000005ad_blk000005b0_Q31_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk000005bc_blk000005bd_blk000005c0_Q31_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk000005c2_blk000005c3_blk000005c5_Q15_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk000005f1_blk00000653_Q15_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk0000091a_blk0000091b_blk0000091e_Q15_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk000009b1_blk000009b2_blk000009cb_Q15_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk000009b1_blk000009b2_blk000009c9_Q15_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk000009b1_blk000009b2_blk000009c7_Q15_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk000009b1_blk000009b2_blk000009c5_Q15_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk000009b1_blk000009b2_blk000009c3_Q15_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk000009b1_blk000009b2_blk000009c1_Q15_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk000009b1_blk000009b2_blk000009bf_Q15_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk000009b1_blk000009b2_blk000009bd_Q15_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk000009b1_blk000009b2_blk000009bb_Q15_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk000009b1_blk000009b2_blk000009b9_Q15_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk000009b1_blk000009b2_blk000009b7_Q15_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk000009b1_blk000009b2_blk000009b5_Q15_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk000009cd_blk000009ce_blk000009e7_Q15_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk000009cd_blk000009ce_blk000009e5_Q15_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk000009cd_blk000009ce_blk000009e3_Q15_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk000009cd_blk000009ce_blk000009e1_Q15_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk000009cd_blk000009ce_blk000009df_Q15_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk000009cd_blk000009ce_blk000009dd_Q15_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk000009cd_blk000009ce_blk000009db_Q15_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk000009cd_blk000009ce_blk000009d9_Q15_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk000009cd_blk000009ce_blk000009d7_Q15_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk000009cd_blk000009ce_blk000009d5_Q15_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk000009cd_blk000009ce_blk000009d3_Q15_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk000009cd_blk000009ce_blk000009d1_Q15_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk000009e9_blk000009ea_blk000009ed_Q15_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000a59_blk00000a5a_blk00000a75_Q15_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000a59_blk00000a5a_blk00000a73_Q15_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000a59_blk00000a5a_blk00000a71_Q15_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000a59_blk00000a5a_blk00000a6f_Q15_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000a59_blk00000a5a_blk00000a6d_Q15_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000a59_blk00000a5a_blk00000a6b_Q15_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000a59_blk00000a5a_blk00000a69_Q15_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000a59_blk00000a5a_blk00000a67_Q15_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000a59_blk00000a5a_blk00000a65_Q15_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000a59_blk00000a5a_blk00000a63_Q15_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000a59_blk00000a5a_blk00000a61_Q15_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000a59_blk00000a5a_blk00000a5f_Q15_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000a59_blk00000a5a_blk00000a5d_Q15_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000a77_blk00000a78_blk00000a93_Q15_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000a77_blk00000a78_blk00000a91_Q15_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000a77_blk00000a78_blk00000a8f_Q15_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000a77_blk00000a78_blk00000a8d_Q15_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000a77_blk00000a78_blk00000a8b_Q15_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000a77_blk00000a78_blk00000a89_Q15_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000a77_blk00000a78_blk00000a87_Q15_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000a77_blk00000a78_blk00000a85_Q15_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000a77_blk00000a78_blk00000a83_Q15_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000a77_blk00000a78_blk00000a81_Q15_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000a77_blk00000a78_blk00000a7f_Q15_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000a77_blk00000a78_blk00000a7d_Q15_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000a77_blk00000a78_blk00000a7b_Q15_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000a95_blk00000a96_blk00000a9b_Q31_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000a95_blk00000a96_blk00000a99_Q31_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000a9d_blk00000a9e_blk00000aa1_Q31_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000aa3_blk00000aa4_blk00000aa7_Q15_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000aa9_blk00000aaa_blk00000aad_Q31_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000aaf_blk00000ab0_blk00000ab5_Q31_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000aaf_blk00000ab0_blk00000ab3_Q31_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000ab7_blk00000ab8_blk00000abd_Q31_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000ab7_blk00000ab8_blk00000abb_Q31_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000abf_blk00000ac0_blk00000acd_Q31_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000abf_blk00000ac0_blk00000acb_Q31_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000abf_blk00000ac0_blk00000ac9_Q31_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000abf_blk00000ac0_blk00000ac7_Q31_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000abf_blk00000ac0_blk00000ac5_Q31_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000abf_blk00000ac0_blk00000ac3_Q31_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000acf_blk00000ad0_blk00000ad5_Q15_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000acf_blk00000ad0_blk00000ad3_Q15_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000b49_blk00000b4a_blk00000b4c_Q15_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000b4e_blk00000b4f_blk00000b51_Q15_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000b53_blk00000b54_blk00000b57_Q15_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000c06_blk00000c07_blk00000c24_Q15_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000c06_blk00000c07_blk00000c22_Q15_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000c06_blk00000c07_blk00000c20_Q15_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000c06_blk00000c07_blk00000c1e_Q15_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000c06_blk00000c07_blk00000c1c_Q15_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000c06_blk00000c07_blk00000c1a_Q15_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000c06_blk00000c07_blk00000c18_Q15_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000c06_blk00000c07_blk00000c16_Q15_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000c06_blk00000c07_blk00000c14_Q15_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000c06_blk00000c07_blk00000c12_Q15_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000c06_blk00000c07_blk00000c10_Q15_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000c06_blk00000c07_blk00000c0e_Q15_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000c06_blk00000c07_blk00000c0c_Q15_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000c06_blk00000c07_blk00000c0a_Q15_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000c26_blk00000c27_blk00000c44_Q15_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000c26_blk00000c27_blk00000c42_Q15_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000c26_blk00000c27_blk00000c40_Q15_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000c26_blk00000c27_blk00000c3e_Q15_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000c26_blk00000c27_blk00000c3c_Q15_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000c26_blk00000c27_blk00000c3a_Q15_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000c26_blk00000c27_blk00000c38_Q15_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000c26_blk00000c27_blk00000c36_Q15_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000c26_blk00000c27_blk00000c34_Q15_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000c26_blk00000c27_blk00000c32_Q15_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000c26_blk00000c27_blk00000c30_Q15_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000c26_blk00000c27_blk00000c2e_Q15_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000c26_blk00000c27_blk00000c2c_Q15_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000c26_blk00000c27_blk00000c2a_Q15_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000c46_blk00000c47_blk00000c64_Q15_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000c46_blk00000c47_blk00000c62_Q15_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000c46_blk00000c47_blk00000c60_Q15_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000c46_blk00000c47_blk00000c5e_Q15_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000c46_blk00000c47_blk00000c5c_Q15_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000c46_blk00000c47_blk00000c5a_Q15_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000c46_blk00000c47_blk00000c58_Q15_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000c46_blk00000c47_blk00000c56_Q15_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000c46_blk00000c47_blk00000c54_Q15_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000c46_blk00000c47_blk00000c52_Q15_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000c46_blk00000c47_blk00000c50_Q15_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000c46_blk00000c47_blk00000c4e_Q15_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000c46_blk00000c47_blk00000c4c_Q15_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000c46_blk00000c47_blk00000c4a_Q15_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000c66_blk00000c67_blk00000c84_Q15_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000c66_blk00000c67_blk00000c82_Q15_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000c66_blk00000c67_blk00000c80_Q15_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000c66_blk00000c67_blk00000c7e_Q15_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000c66_blk00000c67_blk00000c7c_Q15_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000c66_blk00000c67_blk00000c7a_Q15_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000c66_blk00000c67_blk00000c78_Q15_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000c66_blk00000c67_blk00000c76_Q15_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000c66_blk00000c67_blk00000c74_Q15_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000c66_blk00000c67_blk00000c72_Q15_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000c66_blk00000c67_blk00000c70_Q15_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000c66_blk00000c67_blk00000c6e_Q15_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000c66_blk00000c67_blk00000c6c_Q15_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000c66_blk00000c67_blk00000c6a_Q15_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000c86_blk00000c87_blk00000c90_Q15_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000c86_blk00000c87_blk00000c8e_Q15_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000c86_blk00000c87_blk00000c8c_Q15_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000c86_blk00000c87_blk00000c8a_Q15_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000c92_blk00000c93_blk00000c95_Q15_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000cb3_blk00000cd4_Q15_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000cb3_blk00000cd2_Q15_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000cd6_blk00000cd7_blk00000ce4_Q15_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000cd6_blk00000cd7_blk00000ce2_Q15_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000cd6_blk00000cd7_blk00000ce0_Q15_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000cd6_blk00000cd7_blk00000cde_Q15_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000cd6_blk00000cd7_blk00000cdc_Q15_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000cd6_blk00000cd7_blk00000cda_Q15_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000ce6_blk00000ce7_blk00000cea_Q15_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000d58_blk00000d59_blk00000d5b_Q15_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000d91_blk00000d92_blk00000daa_Q15_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000d91_blk00000d92_blk00000da8_Q15_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000d91_blk00000d92_blk00000da6_Q15_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000d91_blk00000d92_blk00000da4_Q15_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000d91_blk00000d92_blk00000da2_Q15_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000d91_blk00000d92_blk00000da0_Q15_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000d91_blk00000d92_blk00000d9e_Q15_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000d91_blk00000d92_blk00000d9c_Q15_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000d91_blk00000d92_blk00000d9a_Q15_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000d91_blk00000d92_blk00000d98_Q15_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000d91_blk00000d92_blk00000d96_Q15_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000d91_blk00000d92_blk00000d94_Q15_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000dac_blk00000dad_blk00000dc5_Q15_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000dac_blk00000dad_blk00000dc3_Q15_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000dac_blk00000dad_blk00000dc1_Q15_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000dac_blk00000dad_blk00000dbf_Q15_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000dac_blk00000dad_blk00000dbd_Q15_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000dac_blk00000dad_blk00000dbb_Q15_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000dac_blk00000dad_blk00000db9_Q15_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000dac_blk00000dad_blk00000db7_Q15_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000dac_blk00000dad_blk00000db5_Q15_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000dac_blk00000dad_blk00000db3_Q15_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000dac_blk00000dad_blk00000db1_Q15_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000dac_blk00000dad_blk00000daf_Q15_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000dc7_blk00000dc8_blk00000de2_Q15_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000dc7_blk00000dc8_blk00000de0_Q15_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000dc7_blk00000dc8_blk00000dde_Q15_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000dc7_blk00000dc8_blk00000ddc_Q15_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000dc7_blk00000dc8_blk00000dda_Q15_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000dc7_blk00000dc8_blk00000dd8_Q15_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000dc7_blk00000dc8_blk00000dd6_Q15_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000dc7_blk00000dc8_blk00000dd4_Q15_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000dc7_blk00000dc8_blk00000dd2_Q15_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000dc7_blk00000dc8_blk00000dd0_Q15_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000dc7_blk00000dc8_blk00000dce_Q15_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000dc7_blk00000dc8_blk00000dcc_Q15_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000dc7_blk00000dc8_blk00000dca_Q15_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000de4_blk00000de5_blk00000dff_Q15_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000de4_blk00000de5_blk00000dfd_Q15_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000de4_blk00000de5_blk00000dfb_Q15_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000de4_blk00000de5_blk00000df9_Q15_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000de4_blk00000de5_blk00000df7_Q15_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000de4_blk00000de5_blk00000df5_Q15_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000de4_blk00000de5_blk00000df3_Q15_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000de4_blk00000de5_blk00000df1_Q15_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000de4_blk00000de5_blk00000def_Q15_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000de4_blk00000de5_blk00000ded_Q15_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000de4_blk00000de5_blk00000deb_Q15_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000de4_blk00000de5_blk00000de9_Q15_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000de4_blk00000de5_blk00000de7_Q15_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000e01_blk00000e02_blk00000e07_Q15_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000e01_blk00000e02_blk00000e05_Q15_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000e09_blk00000e0a_blk00000e0f_Q15_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000e09_blk00000e0a_blk00000e0d_Q15_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000e11_blk00000e12_blk00000e15_Q15_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000e17_blk00000e18_blk00000e1b_Q15_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000e1d_blk00000e1e_blk00000e23_Q15_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000e1d_blk00000e1e_blk00000e21_Q15_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000e25_blk00000e26_blk00000e33_Q15_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000e25_blk00000e26_blk00000e31_Q15_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000e25_blk00000e26_blk00000e2f_Q15_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000e25_blk00000e26_blk00000e2d_Q15_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000e25_blk00000e26_blk00000e2b_Q15_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000e25_blk00000e26_blk00000e29_Q15_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000ea7_blk00000ea8_blk00000eaa_Q15_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000eac_blk00000ead_blk00000eaf_Q15_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000fbf_blk00000fc1_DO_31_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000fbf_blk00000fc1_DO_30_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000fbf_blk00000fc1_DO_29_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000fbf_blk00000fc1_DO_28_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000fbf_blk00000fc1_DO_27_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000fbf_blk00000fc1_DO_26_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000fbf_blk00000fc1_DO_25_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000fbf_blk00000fc1_DO_24_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000fbf_blk00000fc1_DO_23_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000fbf_blk00000fc1_DO_22_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000fbf_blk00000fc1_DOP_3_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000fbf_blk00000fc1_DOP_2_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000fc2_blk00000fc3_blk00000fd0_Q15_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000fc2_blk00000fc3_blk00000fce_Q15_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000fc2_blk00000fc3_blk00000fcc_Q15_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000fc2_blk00000fc3_blk00000fca_Q15_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000fc2_blk00000fc3_blk00000fc8_Q15_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000fc2_blk00000fc3_blk00000fc6_Q15_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000fd8_blk00000fd9_blk00000fdb_Q15_UNCONNECTED : STD_LOGIC; 
  signal NlwRenamedSig_OI_xn_index : STD_LOGIC_VECTOR ( 5 downto 0 ); 
  signal NlwRenamedSig_OI_xk_index : STD_LOGIC_VECTOR ( 5 downto 0 ); 
  signal U0_i_synth_non_floating_point_arch_d_xfft_inst_pe_natural_out : STD_LOGIC_VECTOR ( 23 downto 0 ); 
begin
  xn_index(5) <= NlwRenamedSig_OI_xn_index(5);
  xn_index(4) <= NlwRenamedSig_OI_xn_index(4);
  xn_index(3) <= NlwRenamedSig_OI_xn_index(3);
  xn_index(2) <= NlwRenamedSig_OI_xn_index(2);
  xn_index(1) <= NlwRenamedSig_OI_xn_index(1);
  xn_index(0) <= NlwRenamedSig_OI_xn_index(0);
  xk_index(5) <= NlwRenamedSig_OI_xk_index(5);
  xk_index(4) <= NlwRenamedSig_OI_xk_index(4);
  xk_index(3) <= NlwRenamedSig_OI_xk_index(3);
  xk_index(2) <= NlwRenamedSig_OI_xk_index(2);
  xk_index(1) <= NlwRenamedSig_OI_xk_index(1);
  xk_index(0) <= NlwRenamedSig_OI_xk_index(0);
  xk_re(11) <= U0_i_synth_non_floating_point_arch_d_xfft_inst_pe_natural_out(23);
  xk_re(10) <= U0_i_synth_non_floating_point_arch_d_xfft_inst_pe_natural_out(22);
  xk_re(9) <= U0_i_synth_non_floating_point_arch_d_xfft_inst_pe_natural_out(21);
  xk_re(8) <= U0_i_synth_non_floating_point_arch_d_xfft_inst_pe_natural_out(20);
  xk_re(7) <= U0_i_synth_non_floating_point_arch_d_xfft_inst_pe_natural_out(19);
  xk_re(6) <= U0_i_synth_non_floating_point_arch_d_xfft_inst_pe_natural_out(18);
  xk_re(5) <= U0_i_synth_non_floating_point_arch_d_xfft_inst_pe_natural_out(17);
  xk_re(4) <= U0_i_synth_non_floating_point_arch_d_xfft_inst_pe_natural_out(16);
  xk_re(3) <= U0_i_synth_non_floating_point_arch_d_xfft_inst_pe_natural_out(15);
  xk_re(2) <= U0_i_synth_non_floating_point_arch_d_xfft_inst_pe_natural_out(14);
  xk_re(1) <= U0_i_synth_non_floating_point_arch_d_xfft_inst_pe_natural_out(13);
  xk_re(0) <= U0_i_synth_non_floating_point_arch_d_xfft_inst_pe_natural_out(12);
  xk_im(11) <= U0_i_synth_non_floating_point_arch_d_xfft_inst_pe_natural_out(11);
  xk_im(10) <= U0_i_synth_non_floating_point_arch_d_xfft_inst_pe_natural_out(10);
  xk_im(9) <= U0_i_synth_non_floating_point_arch_d_xfft_inst_pe_natural_out(9);
  xk_im(8) <= U0_i_synth_non_floating_point_arch_d_xfft_inst_pe_natural_out(8);
  xk_im(7) <= U0_i_synth_non_floating_point_arch_d_xfft_inst_pe_natural_out(7);
  xk_im(6) <= U0_i_synth_non_floating_point_arch_d_xfft_inst_pe_natural_out(6);
  xk_im(5) <= U0_i_synth_non_floating_point_arch_d_xfft_inst_pe_natural_out(5);
  xk_im(4) <= U0_i_synth_non_floating_point_arch_d_xfft_inst_pe_natural_out(4);
  xk_im(3) <= U0_i_synth_non_floating_point_arch_d_xfft_inst_pe_natural_out(3);
  xk_im(2) <= U0_i_synth_non_floating_point_arch_d_xfft_inst_pe_natural_out(2);
  xk_im(1) <= U0_i_synth_non_floating_point_arch_d_xfft_inst_pe_natural_out(1);
  xk_im(0) <= U0_i_synth_non_floating_point_arch_d_xfft_inst_pe_natural_out(0);
  rfd <= NlwRenamedSig_OI_U0_i_synth_non_floating_point_arch_d_xfft_inst_FLOW_load_enable;
  busy <= U0_i_synth_non_floating_point_arch_d_xfft_inst_has_bit_reverse_busy_gen_busy_i;
  edone <= NlwRenamedSig_OI_U0_i_synth_non_floating_point_arch_d_xfft_inst_done_int_d;
  done <= U0_i_synth_non_floating_point_arch_d_xfft_inst_DONE;
  dv <= U0_i_synth_non_floating_point_arch_d_xfft_inst_DV;
  cpv <= NlwRenamedSig_OI_cpv;
  rfs <= NlwRenamedSig_OI_rfs;
  blk00000001 : VCC
    port map (
      P => sig000006d1
    );
  blk00000002 : GND
    port map (
      G => sig000008b6
    );
  blk00000003 : LUT3
    generic map(
      INIT => X"AE"
    )
    port map (
      I0 => sig00000042,
      I1 => sig000000a3,
      I2 => sig000000a2,
      O => sig00000014
    );
  blk00000004 : LUT3
    generic map(
      INIT => X"AE"
    )
    port map (
      I0 => sig000000aa,
      I1 => sig00000115,
      I2 => sig00000114,
      O => sig00000018
    );
  blk00000005 : MUXCY
    port map (
      CI => sig000006d1,
      DI => sig000008b6,
      S => sig0000001a,
      O => sig00000019
    );
  blk00000006 : XORCY
    port map (
      CI => sig00000024,
      LI => sig000008b6,
      O => sig00000022
    );
  blk00000007 : MUXCY
    port map (
      CI => sig000006d1,
      DI => sig000008b6,
      S => sig00000025,
      O => sig00000023
    );
  blk00000008 : MUXCY
    port map (
      CI => sig00000023,
      DI => sig000008b6,
      S => sig00000026,
      O => sig00000024
    );
  blk00000009 : LUT6
    generic map(
      INIT => X"9009000000009009"
    )
    port map (
      I0 => sig0000011b,
      I1 => sig000006d1,
      I2 => sig0000011a,
      I3 => sig000008b6,
      I4 => sig00000119,
      I5 => sig000006d1,
      O => sig00000025
    );
  blk0000000a : LUT6
    generic map(
      INIT => X"9009000000009009"
    )
    port map (
      I0 => sig00000118,
      I1 => sig000006d1,
      I2 => sig00000117,
      I3 => sig000006d1,
      I4 => sig00000116,
      I5 => sig000006d1,
      O => sig00000026
    );
  blk0000000b : LUT6
    generic map(
      INIT => X"9009000000009009"
    )
    port map (
      I0 => sig000000c6,
      I1 => sig000006d1,
      I2 => sig000000c7,
      I3 => sig000006d1,
      I4 => sig000000c8,
      I5 => sig000006d1,
      O => sig00000027
    );
  blk0000000c : LUT6
    generic map(
      INIT => X"9009000000009009"
    )
    port map (
      I0 => sig000000c3,
      I1 => sig000006d1,
      I2 => sig000000c4,
      I3 => sig000008b6,
      I4 => sig000000c5,
      I5 => sig000006d1,
      O => sig00000028
    );
  blk0000000d : MUXCY
    port map (
      CI => sig0000002a,
      DI => sig000008b6,
      S => sig00000027,
      O => sig00000029
    );
  blk0000000e : MUXCY
    port map (
      CI => sig000006d1,
      DI => sig000008b6,
      S => sig00000028,
      O => sig0000002a
    );
  blk0000000f : XORCY
    port map (
      CI => sig00000029,
      LI => sig000008b6,
      O => sig00000041
    );
  blk00000010 : LUT6
    generic map(
      INIT => X"9009000000009009"
    )
    port map (
      I0 => sig000000c6,
      I1 => sig000006d1,
      I2 => sig000000c7,
      I3 => sig000006d1,
      I4 => sig000000c8,
      I5 => sig000006d1,
      O => sig0000002b
    );
  blk00000011 : LUT6
    generic map(
      INIT => X"9009000000009009"
    )
    port map (
      I0 => sig000000c3,
      I1 => sig000008b6,
      I2 => sig000000c4,
      I3 => sig000006d1,
      I4 => sig000000c5,
      I5 => sig000006d1,
      O => sig0000002c
    );
  blk00000012 : MUXCY
    port map (
      CI => sig0000002e,
      DI => sig000008b6,
      S => sig0000002b,
      O => sig0000002d
    );
  blk00000013 : MUXCY
    port map (
      CI => sig000006d1,
      DI => sig000008b6,
      S => sig0000002c,
      O => sig0000002e
    );
  blk00000014 : XORCY
    port map (
      CI => sig0000002d,
      LI => sig000008b6,
      O => sig00000040
    );
  blk00000015 : LUT6
    generic map(
      INIT => X"9009000000009009"
    )
    port map (
      I0 => sig000000c6,
      I1 => sig000006d1,
      I2 => sig000000c7,
      I3 => sig000006d1,
      I4 => sig000000c8,
      I5 => sig000006d1,
      O => sig0000002f
    );
  blk00000016 : LUT6
    generic map(
      INIT => X"9009000000009009"
    )
    port map (
      I0 => sig000000c3,
      I1 => sig000006d1,
      I2 => sig000000c4,
      I3 => sig000006d1,
      I4 => sig000000c5,
      I5 => sig000006d1,
      O => sig00000030
    );
  blk00000017 : MUXCY
    port map (
      CI => sig00000032,
      DI => sig000008b6,
      S => sig0000002f,
      O => sig00000031
    );
  blk00000018 : MUXCY
    port map (
      CI => sig000006d1,
      DI => sig000008b6,
      S => sig00000030,
      O => sig00000032
    );
  blk00000019 : XORCY
    port map (
      CI => sig00000031,
      LI => sig000008b6,
      O => sig0000003f
    );
  blk0000001a : FDR
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      D => sig00000002,
      R => sig000008b6,
      Q => sig00000061
    );
  blk0000001b : FDR
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      D => sig00000004,
      R => sig000008b6,
      Q => sig00000062
    );
  blk0000001c : FDR
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      D => sig00000006,
      R => sig000008b6,
      Q => NlwRenamedSig_OI_cpv
    );
  blk0000001d : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => sig0000011b,
      Q => sig00000051
    );
  blk0000001e : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => sig0000011a,
      Q => sig00000050
    );
  blk0000001f : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => sig00000119,
      Q => sig0000004f
    );
  blk00000020 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => sig00000118,
      Q => sig0000004e
    );
  blk00000021 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => sig00000117,
      Q => sig0000004d
    );
  blk00000022 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => sig00000116,
      Q => sig0000004c
    );
  blk00000023 : FDR
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      D => sig00000007,
      R => sig000008b6,
      Q => sig000000a0
    );
  blk00000024 : FDR
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      D => sig00000008,
      R => sig000008b6,
      Q => sig0000009f
    );
  blk00000025 : FDR
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      D => sig00000009,
      R => sig000008b6,
      Q => sig0000009e
    );
  blk00000026 : FDR
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      D => sig0000000a,
      R => sig000008b6,
      Q => sig0000009d
    );
  blk00000027 : FDR
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      D => sig0000000b,
      R => sig000008b6,
      Q => sig0000009c
    );
  blk00000028 : FDR
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      D => sig0000000c,
      R => sig000008b6,
      Q => sig0000009b
    );
  blk00000029 : FDR
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      D => sig0000000d,
      R => sig000008b6,
      Q => sig00000093
    );
  blk0000002a : FDR
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      D => sig0000000e,
      R => sig000008b6,
      Q => sig00000094
    );
  blk0000002b : FDR
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      D => sig0000000f,
      R => sig000008b6,
      Q => sig00000095
    );
  blk0000002c : FDR
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      D => sig00000010,
      R => sig000008b6,
      Q => sig00000096
    );
  blk0000002d : FDR
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      D => sig00000011,
      R => sig000008b6,
      Q => sig00000097
    );
  blk0000002e : FDR
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      D => sig00000012,
      R => sig000008b6,
      Q => sig00000098
    );
  blk0000002f : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => sig00000014,
      R => sig000008b6,
      Q => sig000000a3
    );
  blk00000030 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => sig00000046,
      Q => sig0000009a
    );
  blk00000031 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => sig00000045,
      Q => sig00000099
    );
  blk00000032 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => sig0000011d,
      Q => sig00000015
    );
  blk00000033 : FDR
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      D => sig00000016,
      R => sig000008b6,
      Q => sig00000112
    );
  blk00000034 : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => sig00000018,
      R => sig000008b6,
      Q => sig00000115
    );
  blk00000035 : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => sig00000017,
      D => sig00000022,
      R => sig000008b6,
      Q => sig00000021
    );
  blk00000036 : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => sig00000017,
      D => sig00000021,
      R => sig000008b6,
      Q => sig00000114
    );
  blk00000037 : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => sig0000007a,
      R => sig00000044,
      Q => U0_i_synth_non_floating_point_arch_d_xfft_inst_pe_natural_out(23)
    );
  blk00000038 : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => sig00000079,
      R => sig00000044,
      Q => U0_i_synth_non_floating_point_arch_d_xfft_inst_pe_natural_out(22)
    );
  blk00000039 : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => sig00000078,
      R => sig00000044,
      Q => U0_i_synth_non_floating_point_arch_d_xfft_inst_pe_natural_out(21)
    );
  blk0000003a : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => sig00000077,
      R => sig00000044,
      Q => U0_i_synth_non_floating_point_arch_d_xfft_inst_pe_natural_out(20)
    );
  blk0000003b : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => sig00000076,
      R => sig00000044,
      Q => U0_i_synth_non_floating_point_arch_d_xfft_inst_pe_natural_out(19)
    );
  blk0000003c : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => sig00000075,
      R => sig00000044,
      Q => U0_i_synth_non_floating_point_arch_d_xfft_inst_pe_natural_out(18)
    );
  blk0000003d : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => sig00000074,
      R => sig00000044,
      Q => U0_i_synth_non_floating_point_arch_d_xfft_inst_pe_natural_out(17)
    );
  blk0000003e : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => sig00000073,
      R => sig00000044,
      Q => U0_i_synth_non_floating_point_arch_d_xfft_inst_pe_natural_out(16)
    );
  blk0000003f : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => sig00000072,
      R => sig00000044,
      Q => U0_i_synth_non_floating_point_arch_d_xfft_inst_pe_natural_out(15)
    );
  blk00000040 : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => sig00000071,
      R => sig00000044,
      Q => U0_i_synth_non_floating_point_arch_d_xfft_inst_pe_natural_out(14)
    );
  blk00000041 : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => sig00000070,
      R => sig00000044,
      Q => U0_i_synth_non_floating_point_arch_d_xfft_inst_pe_natural_out(13)
    );
  blk00000042 : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => sig0000006f,
      R => sig00000044,
      Q => U0_i_synth_non_floating_point_arch_d_xfft_inst_pe_natural_out(12)
    );
  blk00000043 : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => sig0000006e,
      R => sig00000044,
      Q => U0_i_synth_non_floating_point_arch_d_xfft_inst_pe_natural_out(11)
    );
  blk00000044 : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => sig0000006d,
      R => sig00000044,
      Q => U0_i_synth_non_floating_point_arch_d_xfft_inst_pe_natural_out(10)
    );
  blk00000045 : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => sig0000006c,
      R => sig00000044,
      Q => U0_i_synth_non_floating_point_arch_d_xfft_inst_pe_natural_out(9)
    );
  blk00000046 : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => sig0000006b,
      R => sig00000044,
      Q => U0_i_synth_non_floating_point_arch_d_xfft_inst_pe_natural_out(8)
    );
  blk00000047 : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => sig0000006a,
      R => sig00000044,
      Q => U0_i_synth_non_floating_point_arch_d_xfft_inst_pe_natural_out(7)
    );
  blk00000048 : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => sig00000069,
      R => sig00000044,
      Q => U0_i_synth_non_floating_point_arch_d_xfft_inst_pe_natural_out(6)
    );
  blk00000049 : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => sig00000068,
      R => sig00000044,
      Q => U0_i_synth_non_floating_point_arch_d_xfft_inst_pe_natural_out(5)
    );
  blk0000004a : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => sig00000067,
      R => sig00000044,
      Q => U0_i_synth_non_floating_point_arch_d_xfft_inst_pe_natural_out(4)
    );
  blk0000004b : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => sig00000066,
      R => sig00000044,
      Q => U0_i_synth_non_floating_point_arch_d_xfft_inst_pe_natural_out(3)
    );
  blk0000004c : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => sig00000065,
      R => sig00000044,
      Q => U0_i_synth_non_floating_point_arch_d_xfft_inst_pe_natural_out(2)
    );
  blk0000004d : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => sig00000064,
      R => sig00000044,
      Q => U0_i_synth_non_floating_point_arch_d_xfft_inst_pe_natural_out(1)
    );
  blk0000004e : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => sig00000063,
      R => sig00000044,
      Q => U0_i_synth_non_floating_point_arch_d_xfft_inst_pe_natural_out(0)
    );
  blk0000004f : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => sig00000047,
      R => sig000008b6,
      Q => sig00000048
    );
  blk00000050 : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => sig00000049,
      R => sig000008b6,
      Q => U0_i_synth_non_floating_point_arch_d_xfft_inst_DV
    );
  blk00000051 : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => NlwRenamedSig_OI_U0_i_synth_non_floating_point_arch_d_xfft_inst_done_int_d,
      R => sig000008b6,
      Q => U0_i_synth_non_floating_point_arch_d_xfft_inst_DONE
    );
  blk00000052 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => sig00000038,
      Q => sig0000005d
    );
  blk00000053 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => sig00000037,
      Q => sig0000005c
    );
  blk00000054 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => sig00000036,
      Q => sig0000005b
    );
  blk00000055 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => sig00000035,
      Q => sig0000005a
    );
  blk00000056 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => sig00000034,
      Q => sig00000059
    );
  blk00000057 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => sig00000033,
      Q => sig00000058
    );
  blk00000058 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => sig0000003e,
      Q => sig00000057
    );
  blk00000059 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => sig0000003d,
      Q => sig00000056
    );
  blk0000005a : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => sig0000003c,
      Q => sig00000055
    );
  blk0000005b : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => sig0000003b,
      Q => sig00000054
    );
  blk0000005c : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => sig0000003a,
      Q => sig00000053
    );
  blk0000005d : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => sig00000039,
      Q => sig00000052
    );
  blk0000005e : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => sig00000061,
      R => sig000008b6,
      Q => sig00000049
    );
  blk0000005f : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => sig00000062,
      R => sig000008b6,
      Q => NlwRenamedSig_OI_U0_i_synth_non_floating_point_arch_d_xfft_inst_done_int_d
    );
  blk00000060 : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => sig00000114,
      R => sig000008b6,
      Q => sig0000004a
    );
  blk00000061 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => sig0000003f,
      Q => sig0000005e
    );
  blk00000062 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => sig00000040,
      Q => sig0000005f
    );
  blk00000063 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => sig00000041,
      Q => sig00000060
    );
  blk00000064 : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => sig000000aa,
      R => sig000008b6,
      Q => sig0000004b
    );
  blk0000009d : LUT6
    generic map(
      INIT => X"9009000000009009"
    )
    port map (
      I0 => sig000006d1,
      I1 => NlwRenamedSig_OI_xn_index(3),
      I2 => sig000006d1,
      I3 => NlwRenamedSig_OI_xn_index(4),
      I4 => sig000008b6,
      I5 => NlwRenamedSig_OI_xn_index(5),
      O => sig00000142
    );
  blk0000009e : LUT6
    generic map(
      INIT => X"9009000000009009"
    )
    port map (
      I0 => sig000006d1,
      I1 => NlwRenamedSig_OI_xn_index(0),
      I2 => sig000006d1,
      I3 => NlwRenamedSig_OI_xn_index(1),
      I4 => sig000006d1,
      I5 => NlwRenamedSig_OI_xn_index(2),
      O => sig00000143
    );
  blk0000009f : MUXCY
    port map (
      CI => sig00000145,
      DI => sig000008b6,
      S => sig00000142,
      O => sig00000144
    );
  blk000000a0 : MUXCY
    port map (
      CI => sig000006d1,
      DI => sig000008b6,
      S => sig00000143,
      O => sig00000145
    );
  blk000000a1 : XORCY
    port map (
      CI => sig00000144,
      LI => sig000008b6,
      O => sig0000017d
    );
  blk000000a2 : LUT6
    generic map(
      INIT => X"9009000000009009"
    )
    port map (
      I0 => NlwRenamedSig_OI_xn_index(3),
      I1 => sig000006d1,
      I2 => NlwRenamedSig_OI_xn_index(4),
      I3 => sig000006d1,
      I4 => NlwRenamedSig_OI_xn_index(5),
      I5 => sig000006d1,
      O => sig00000146
    );
  blk000000a3 : LUT6
    generic map(
      INIT => X"9009000000009009"
    )
    port map (
      I0 => NlwRenamedSig_OI_xn_index(0),
      I1 => sig000006d1,
      I2 => NlwRenamedSig_OI_xn_index(1),
      I3 => sig000008b6,
      I4 => NlwRenamedSig_OI_xn_index(2),
      I5 => sig000006d1,
      O => sig00000147
    );
  blk000000a4 : MUXCY
    port map (
      CI => sig00000149,
      DI => sig000008b6,
      S => sig00000146,
      O => sig00000148
    );
  blk000000a5 : MUXCY
    port map (
      CI => sig000006d1,
      DI => sig000008b6,
      S => sig00000147,
      O => sig00000149
    );
  blk000000a6 : XORCY
    port map (
      CI => sig00000148,
      LI => sig000008b6,
      O => sig0000017c
    );
  blk000000a7 : LUT6
    generic map(
      INIT => X"9009000000009009"
    )
    port map (
      I0 => sig00000195,
      I1 => sig000006d1,
      I2 => sig00000196,
      I3 => sig000006d1,
      I4 => sig00000197,
      I5 => sig000006d1,
      O => sig0000014a
    );
  blk000000a8 : LUT6
    generic map(
      INIT => X"9009000000009009"
    )
    port map (
      I0 => sig00000192,
      I1 => sig000006d1,
      I2 => sig00000193,
      I3 => sig000008b6,
      I4 => sig00000194,
      I5 => sig000006d1,
      O => sig0000014b
    );
  blk000000a9 : MUXCY
    port map (
      CI => sig0000014d,
      DI => sig000008b6,
      S => sig0000014a,
      O => sig0000014c
    );
  blk000000aa : MUXCY
    port map (
      CI => sig000006d1,
      DI => sig000008b6,
      S => sig0000014b,
      O => sig0000014d
    );
  blk000000ab : XORCY
    port map (
      CI => sig0000014c,
      LI => sig000008b6,
      O => sig0000017a
    );
  blk000000ac : LUT6
    generic map(
      INIT => X"9009000000009009"
    )
    port map (
      I0 => sig00000121,
      I1 => sig000006d1,
      I2 => sig00000122,
      I3 => sig000006d1,
      I4 => sig00000123,
      I5 => sig000006d1,
      O => sig0000014e
    );
  blk000000ad : LUT6
    generic map(
      INIT => X"9009000000009009"
    )
    port map (
      I0 => sig0000011e,
      I1 => sig000006d1,
      I2 => sig0000011f,
      I3 => sig000008b6,
      I4 => sig00000120,
      I5 => sig000006d1,
      O => sig0000014f
    );
  blk000000ae : MUXCY
    port map (
      CI => sig00000151,
      DI => sig000008b6,
      S => sig0000014e,
      O => sig00000150
    );
  blk000000af : MUXCY
    port map (
      CI => sig000006d1,
      DI => sig000008b6,
      S => sig0000014f,
      O => sig00000151
    );
  blk000000b0 : XORCY
    port map (
      CI => sig00000150,
      LI => sig000008b6,
      O => sig00000175
    );
  blk000000b1 : LUT6
    generic map(
      INIT => X"9009000000009009"
    )
    port map (
      I0 => sig00000121,
      I1 => sig000006d1,
      I2 => sig00000122,
      I3 => sig000006d1,
      I4 => sig00000123,
      I5 => sig000006d1,
      O => sig00000152
    );
  blk000000b2 : LUT6
    generic map(
      INIT => X"9009000000009009"
    )
    port map (
      I0 => sig0000011e,
      I1 => sig000008b6,
      I2 => sig0000011f,
      I3 => sig000006d1,
      I4 => sig00000120,
      I5 => sig000006d1,
      O => sig00000153
    );
  blk000000b3 : MUXCY
    port map (
      CI => sig00000155,
      DI => sig000008b6,
      S => sig00000152,
      O => sig00000154
    );
  blk000000b4 : MUXCY
    port map (
      CI => sig000006d1,
      DI => sig000008b6,
      S => sig00000153,
      O => sig00000155
    );
  blk000000b5 : XORCY
    port map (
      CI => sig00000154,
      LI => sig000008b6,
      O => sig00000174
    );
  blk000000b6 : LUT6
    generic map(
      INIT => X"9009000000009009"
    )
    port map (
      I0 => sig00000121,
      I1 => sig000006d1,
      I2 => sig00000122,
      I3 => sig000006d1,
      I4 => sig00000123,
      I5 => sig000006d1,
      O => sig00000156
    );
  blk000000b7 : LUT6
    generic map(
      INIT => X"9009000000009009"
    )
    port map (
      I0 => sig0000011e,
      I1 => sig000006d1,
      I2 => sig0000011f,
      I3 => sig000006d1,
      I4 => sig00000120,
      I5 => sig000006d1,
      O => sig00000157
    );
  blk000000b8 : MUXCY
    port map (
      CI => sig00000159,
      DI => sig000008b6,
      S => sig00000156,
      O => sig00000158
    );
  blk000000b9 : MUXCY
    port map (
      CI => sig000006d1,
      DI => sig000008b6,
      S => sig00000157,
      O => sig00000159
    );
  blk000000ba : XORCY
    port map (
      CI => sig00000158,
      LI => sig000008b6,
      O => sig00000173
    );
  blk000000bb : LUT6
    generic map(
      INIT => X"9009000000009009"
    )
    port map (
      I0 => NlwRenamedSig_OI_xn_index(3),
      I1 => sig000006d1,
      I2 => NlwRenamedSig_OI_xn_index(4),
      I3 => sig000006d1,
      I4 => NlwRenamedSig_OI_xn_index(5),
      I5 => sig000006d1,
      O => sig0000015a
    );
  blk000000bc : LUT6
    generic map(
      INIT => X"9009000000009009"
    )
    port map (
      I0 => NlwRenamedSig_OI_xn_index(0),
      I1 => sig000006d1,
      I2 => NlwRenamedSig_OI_xn_index(1),
      I3 => sig000008b6,
      I4 => NlwRenamedSig_OI_xn_index(2),
      I5 => sig000006d1,
      O => sig0000015b
    );
  blk000000bd : MUXCY
    port map (
      CI => sig0000015d,
      DI => sig000008b6,
      S => sig0000015a,
      O => sig0000015c
    );
  blk000000be : MUXCY
    port map (
      CI => sig000006d1,
      DI => sig000008b6,
      S => sig0000015b,
      O => sig0000015d
    );
  blk000000bf : XORCY
    port map (
      CI => sig0000015c,
      LI => sig000008b6,
      O => sig0000015e
    );
  blk000000c0 : MUXCY
    port map (
      CI => sig000006d1,
      DI => sig000008b6,
      S => sig00000166,
      O => sig00000167
    );
  blk000000c1 : XORCY
    port map (
      CI => sig0000016d,
      LI => sig000008b6,
      O => sig0000016b
    );
  blk000000c2 : MUXCY
    port map (
      CI => sig000006d1,
      DI => sig000008b6,
      S => sig00000176,
      O => sig0000016c
    );
  blk000000c3 : MUXCY
    port map (
      CI => sig00000179,
      DI => sig000008b6,
      S => sig0000016f,
      O => sig0000016d
    );
  blk000000c4 : MUXCY
    port map (
      CI => sig0000017b,
      DI => sig0000018e,
      S => sig00000171,
      O => sig00000177
    );
  blk000000c5 : MUXCY
    port map (
      CI => sig00000177,
      DI => NlwRenamedSig_OI_rfs,
      S => sig00000178,
      O => sig00000179
    );
  blk000000c6 : MUXCY
    port map (
      CI => sig0000016c,
      DI => sig00000198,
      S => sig00000172,
      O => sig0000017b
    );
  blk000000c7 : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => sig00000186,
      D => sig0000015f,
      R => sig000008b6,
      Q => sig00000198
    );
  blk000000c8 : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => sig00000186,
      D => sig0000015e,
      R => sig000008b6,
      Q => sig0000015f
    );
  blk000000c9 : FDSE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => sig0000016b,
      S => sig000008b6,
      Q => NlwRenamedSig_OI_rfs
    );
  blk000000ca : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => sig0000017a,
      Q => sig0000018d
    );
  blk000000cb : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => sig00000173,
      Q => sig00000187
    );
  blk000000cc : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => sig00000174,
      Q => sig00000188
    );
  blk000000cd : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => sig00000175,
      Q => sig00000189
    );
  blk000000ce : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => sig0000017c,
      Q => sig0000018e
    );
  blk000000cf : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => sig0000017d,
      Q => sig0000011d
    );
  blk000000d0 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => sig00000168,
      D => sig000001a4,
      Q => sig00000129
    );
  blk000000d1 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => sig00000168,
      D => sig000001a3,
      Q => sig00000128
    );
  blk000000d2 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => sig00000168,
      D => sig000001a2,
      Q => sig00000127
    );
  blk000000d3 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => sig00000168,
      D => sig000001a1,
      Q => sig00000126
    );
  blk000000d4 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => sig00000168,
      D => sig000001a0,
      Q => sig00000125
    );
  blk000000d5 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => sig00000168,
      D => sig0000019f,
      Q => sig00000124
    );
  blk000000d6 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => sig00000168,
      D => sig0000018a,
      Q => sig0000011c
    );
  blk000000d7 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => sig00000198,
      Q => sig0000018c
    );
  blk000000d8 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => sig00000170,
      Q => NlwRenamedSig_OI_U0_i_synth_non_floating_point_arch_d_xfft_inst_FLOW_load_enable
    );
  blk000000d9 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => sig00000168,
      D => sig00000183,
      Q => sig00000123
    );
  blk000000da : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => sig00000168,
      D => sig00000182,
      Q => sig00000122
    );
  blk000000db : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => sig00000168,
      D => sig00000181,
      Q => sig00000121
    );
  blk000000dc : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => sig00000168,
      D => sig00000180,
      Q => sig00000120
    );
  blk000000dd : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => sig00000168,
      D => sig0000017f,
      Q => sig0000011f
    );
  blk000000de : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => sig00000168,
      D => sig0000017e,
      Q => sig0000011e
    );
  blk000000df : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => sig00000184,
      Q => sig0000018b
    );
  blk000000e0 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => sig0000016e,
      Q => sig0000018f
    );
  blk000000e1 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => sig00000169,
      D => cp_len(5),
      Q => sig0000019e
    );
  blk000000e2 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => sig00000169,
      D => cp_len(4),
      Q => sig0000019d
    );
  blk000000e3 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => sig00000169,
      D => cp_len(3),
      Q => sig0000019c
    );
  blk000000e4 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => sig00000169,
      D => cp_len(2),
      Q => sig0000019b
    );
  blk000000e5 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => sig00000169,
      D => cp_len(1),
      Q => sig0000019a
    );
  blk000000e6 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => sig00000169,
      D => cp_len(0),
      Q => sig00000199
    );
  blk000000e7 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => sig0000016a,
      D => scale_sch(5),
      Q => sig000001a4
    );
  blk000000e8 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => sig0000016a,
      D => scale_sch(4),
      Q => sig000001a3
    );
  blk000000e9 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => sig0000016a,
      D => scale_sch(3),
      Q => sig000001a2
    );
  blk000000ea : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => sig0000016a,
      D => scale_sch(2),
      Q => sig000001a1
    );
  blk000000eb : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => sig0000016a,
      D => scale_sch(1),
      Q => sig000001a0
    );
  blk000000ec : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => sig0000016a,
      D => scale_sch(0),
      Q => sig0000019f
    );
  blk00000132 : LUT6
    generic map(
      INIT => X"9009000000009009"
    )
    port map (
      I0 => sig00000123,
      I1 => sig000006d1,
      I2 => sig000008b6,
      I3 => sig000008b6,
      I4 => sig000008b6,
      I5 => sig000008b6,
      O => sig000001a5
    );
  blk00000133 : LUT6
    generic map(
      INIT => X"9009000000009009"
    )
    port map (
      I0 => sig00000120,
      I1 => sig000006d1,
      I2 => sig00000121,
      I3 => sig000006d1,
      I4 => sig00000122,
      I5 => sig000006d1,
      O => sig000001a6
    );
  blk00000134 : LUT6
    generic map(
      INIT => X"9009000000009009"
    )
    port map (
      I0 => sig00000198,
      I1 => sig000006d1,
      I2 => sig0000011e,
      I3 => sig000006d1,
      I4 => sig0000011f,
      I5 => sig000008b6,
      O => sig000001a7
    );
  blk00000135 : MUXCY
    port map (
      CI => sig000001a9,
      DI => sig000008b6,
      S => sig000001a5,
      O => sig000001a8
    );
  blk00000136 : MUXCY
    port map (
      CI => sig000001aa,
      DI => sig000008b6,
      S => sig000001a6,
      O => sig000001a9
    );
  blk00000137 : MUXCY
    port map (
      CI => sig000006d1,
      DI => sig000008b6,
      S => sig000001a7,
      O => sig000001aa
    );
  blk00000138 : XORCY
    port map (
      CI => sig000001a8,
      LI => sig000008b6,
      O => sig000001ba
    );
  blk00000139 : LUT6
    generic map(
      INIT => X"9009000000009009"
    )
    port map (
      I0 => sig00000123,
      I1 => sig000006d1,
      I2 => sig000008b6,
      I3 => sig000008b6,
      I4 => sig000008b6,
      I5 => sig000008b6,
      O => sig000001ab
    );
  blk0000013a : LUT6
    generic map(
      INIT => X"9009000000009009"
    )
    port map (
      I0 => sig00000120,
      I1 => sig000006d1,
      I2 => sig00000121,
      I3 => sig000006d1,
      I4 => sig00000122,
      I5 => sig000006d1,
      O => sig000001ac
    );
  blk0000013b : LUT6
    generic map(
      INIT => X"9009000000009009"
    )
    port map (
      I0 => sig00000198,
      I1 => sig000006d1,
      I2 => sig0000011e,
      I3 => sig000008b6,
      I4 => sig0000011f,
      I5 => sig000006d1,
      O => sig000001ad
    );
  blk0000013c : MUXCY
    port map (
      CI => sig000001ae,
      DI => sig000008b6,
      S => sig000001ab,
      O => sig000001bb
    );
  blk0000013d : MUXCY
    port map (
      CI => sig000001af,
      DI => sig000008b6,
      S => sig000001ac,
      O => sig000001ae
    );
  blk0000013e : MUXCY
    port map (
      CI => sig000006d1,
      DI => sig000008b6,
      S => sig000001ad,
      O => sig000001af
    );
  blk0000013f : LUT6
    generic map(
      INIT => X"9009000000009009"
    )
    port map (
      I0 => sig00000195,
      I1 => sig000006d1,
      I2 => sig00000196,
      I3 => sig000006d1,
      I4 => sig00000197,
      I5 => sig000006d1,
      O => sig000001b0
    );
  blk00000140 : LUT6
    generic map(
      INIT => X"9009000000009009"
    )
    port map (
      I0 => sig00000192,
      I1 => sig000006d1,
      I2 => sig00000193,
      I3 => sig000008b6,
      I4 => sig00000194,
      I5 => sig000006d1,
      O => sig000001b1
    );
  blk00000141 : MUXCY
    port map (
      CI => sig000001b3,
      DI => sig000008b6,
      S => sig000001b0,
      O => sig000001b2
    );
  blk00000142 : MUXCY
    port map (
      CI => sig000006d1,
      DI => sig000008b6,
      S => sig000001b1,
      O => sig000001b3
    );
  blk00000143 : XORCY
    port map (
      CI => sig000001b2,
      LI => sig000008b6,
      O => sig000001c5
    );
  blk00000144 : XORCY
    port map (
      CI => sig000001b7,
      LI => sig000008b6,
      O => sig000001b4
    );
  blk00000145 : MUXCY
    port map (
      CI => sig000001bb,
      DI => sig000001bc,
      S => sig000001b6,
      O => sig000001b5
    );
  blk00000146 : MUXCY
    port map (
      CI => sig000001b5,
      DI => sig000001bd,
      S => sig000001b8,
      O => sig000001b7
    );
  blk00000147 : MUXCY
    port map (
      CI => sig000006d1,
      DI => sig000008b6,
      S => sig000001be,
      O => sig000001b9
    );
  blk00000148 : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => sig00000185,
      D => sig000001ba,
      R => sig000008b6,
      Q => sig000001bc
    );
  blk00000149 : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => sig00000185,
      D => sig000001c5,
      R => sig000008b6,
      Q => sig000001bd
    );
  blk0000014a : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => sig00000185,
      D => sig000001b4,
      R => sig000008b6,
      Q => sig00000191
    );
  blk00000162 : LUT6
    generic map(
      INIT => X"9009000000009009"
    )
    port map (
      I0 => sig000000c8,
      I1 => sig000006d1,
      I2 => sig000008b6,
      I3 => sig000008b6,
      I4 => sig000008b6,
      I5 => sig000008b6,
      O => sig000001c6
    );
  blk00000163 : LUT6
    generic map(
      INIT => X"9009000000009009"
    )
    port map (
      I0 => sig000000c5,
      I1 => sig000006d1,
      I2 => sig000000c6,
      I3 => sig000006d1,
      I4 => sig000000c7,
      I5 => sig000006d1,
      O => sig000001c7
    );
  blk00000164 : LUT6
    generic map(
      INIT => X"9009000000009009"
    )
    port map (
      I0 => sig00000043,
      I1 => sig000006d1,
      I2 => sig000000c3,
      I3 => sig000006d1,
      I4 => sig000000c4,
      I5 => sig000008b6,
      O => sig000001c8
    );
  blk00000165 : MUXCY
    port map (
      CI => sig000001ca,
      DI => sig000008b6,
      S => sig000001c6,
      O => sig000001c9
    );
  blk00000166 : MUXCY
    port map (
      CI => sig000001cb,
      DI => sig000008b6,
      S => sig000001c7,
      O => sig000001ca
    );
  blk00000167 : MUXCY
    port map (
      CI => sig000006d1,
      DI => sig000008b6,
      S => sig000001c8,
      O => sig000001cb
    );
  blk00000168 : XORCY
    port map (
      CI => sig000001c9,
      LI => sig000008b6,
      O => sig000001db
    );
  blk00000169 : LUT6
    generic map(
      INIT => X"9009000000009009"
    )
    port map (
      I0 => sig000000c8,
      I1 => sig000006d1,
      I2 => sig000008b6,
      I3 => sig000008b6,
      I4 => sig000008b6,
      I5 => sig000008b6,
      O => sig000001cc
    );
  blk0000016a : LUT6
    generic map(
      INIT => X"9009000000009009"
    )
    port map (
      I0 => sig000000c5,
      I1 => sig000006d1,
      I2 => sig000000c6,
      I3 => sig000006d1,
      I4 => sig000000c7,
      I5 => sig000006d1,
      O => sig000001cd
    );
  blk0000016b : LUT6
    generic map(
      INIT => X"9009000000009009"
    )
    port map (
      I0 => sig00000043,
      I1 => sig000006d1,
      I2 => sig000000c3,
      I3 => sig000008b6,
      I4 => sig000000c4,
      I5 => sig000006d1,
      O => sig000001ce
    );
  blk0000016c : MUXCY
    port map (
      CI => sig000001cf,
      DI => sig000008b6,
      S => sig000001cc,
      O => sig000001dc
    );
  blk0000016d : MUXCY
    port map (
      CI => sig000001d0,
      DI => sig000008b6,
      S => sig000001cd,
      O => sig000001cf
    );
  blk0000016e : MUXCY
    port map (
      CI => sig000006d1,
      DI => sig000008b6,
      S => sig000001ce,
      O => sig000001d0
    );
  blk0000016f : LUT6
    generic map(
      INIT => X"9009000000009009"
    )
    port map (
      I0 => sig000000a7,
      I1 => sig000006d1,
      I2 => sig000000a8,
      I3 => sig000006d1,
      I4 => sig000000a9,
      I5 => sig000006d1,
      O => sig000001d1
    );
  blk00000170 : LUT6
    generic map(
      INIT => X"9009000000009009"
    )
    port map (
      I0 => sig000000a4,
      I1 => sig000006d1,
      I2 => sig000000a5,
      I3 => sig000008b6,
      I4 => sig000000a6,
      I5 => sig000006d1,
      O => sig000001d2
    );
  blk00000171 : MUXCY
    port map (
      CI => sig000001d4,
      DI => sig000008b6,
      S => sig000001d1,
      O => sig000001d3
    );
  blk00000172 : MUXCY
    port map (
      CI => sig000006d1,
      DI => sig000008b6,
      S => sig000001d2,
      O => sig000001d4
    );
  blk00000173 : XORCY
    port map (
      CI => sig000001d3,
      LI => sig000008b6,
      O => sig000001e6
    );
  blk00000174 : XORCY
    port map (
      CI => sig000001d8,
      LI => sig000008b6,
      O => sig000001d5
    );
  blk00000175 : MUXCY
    port map (
      CI => sig000001dc,
      DI => sig000001dd,
      S => sig000001d7,
      O => sig000001d6
    );
  blk00000176 : MUXCY
    port map (
      CI => sig000001d6,
      DI => sig000001de,
      S => sig000001d9,
      O => sig000001d8
    );
  blk00000177 : MUXCY
    port map (
      CI => sig000006d1,
      DI => sig000008b6,
      S => sig000001df,
      O => sig000001da
    );
  blk00000178 : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => sig00000013,
      D => sig000001db,
      R => sig000008b6,
      Q => sig000001dd
    );
  blk00000179 : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => sig00000013,
      D => sig000001e6,
      R => sig000008b6,
      Q => sig000001de
    );
  blk0000017a : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => sig00000013,
      D => sig000001d5,
      R => sig000008b6,
      Q => sig000000a2
    );
  blk0000019b : FDR
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      D => sig000001e8,
      R => sig000008b6,
      Q => sig000000ee
    );
  blk0000019c : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => sig000001ea,
      D => sig00000124,
      Q => sig00000253
    );
  blk0000019d : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => sig000001ea,
      D => sig00000125,
      Q => sig00000254
    );
  blk0000019e : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => sig000001ea,
      D => sig00000126,
      Q => sig00000255
    );
  blk0000019f : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => sig000001ea,
      D => sig00000127,
      Q => sig00000256
    );
  blk000001a0 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => sig000001ea,
      D => sig00000128,
      Q => sig00000257
    );
  blk000001a1 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => sig000001ea,
      D => sig00000129,
      Q => sig00000258
    );
  blk000001a2 : FD
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      D => sig000001e9,
      Q => sig0000025a
    );
  blk000001a3 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => sig000001ea,
      D => sig0000025a,
      Q => sig000001eb
    );
  blk000001a4 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => sig000001ea,
      D => sig00000123,
      Q => sig00000260
    );
  blk000001a5 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => sig000001ea,
      D => sig00000122,
      Q => sig0000025f
    );
  blk000001a6 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => sig000001ea,
      D => sig00000121,
      Q => sig0000025e
    );
  blk000001a7 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => sig000001ea,
      D => sig00000120,
      Q => sig0000025d
    );
  blk000001a8 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => sig000001ea,
      D => sig0000011f,
      Q => sig0000025c
    );
  blk000001a9 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => sig000001ea,
      D => sig0000011e,
      Q => sig0000025b
    );
  blk000001c1 : LUT6
    generic map(
      INIT => X"9009000000009009"
    )
    port map (
      I0 => sig00000286,
      I1 => sig000006d1,
      I2 => sig00000287,
      I3 => sig000008b6,
      I4 => sig00000288,
      I5 => sig000008b6,
      O => sig00000289
    );
  blk000001c2 : LUT6
    generic map(
      INIT => X"9009000000009009"
    )
    port map (
      I0 => sig00000283,
      I1 => sig000008b6,
      I2 => sig00000284,
      I3 => sig000006d1,
      I4 => sig00000285,
      I5 => sig000006d1,
      O => sig0000028a
    );
  blk000001c3 : MUXCY
    port map (
      CI => sig0000028b,
      DI => sig000008b6,
      S => sig00000289,
      O => sig0000029c
    );
  blk000001c4 : MUXCY
    port map (
      CI => sig000006d1,
      DI => sig000008b6,
      S => sig0000028a,
      O => sig0000028b
    );
  blk000001c5 : LUT6
    generic map(
      INIT => X"9009000000009009"
    )
    port map (
      I0 => sig00000286,
      I1 => sig000006d1,
      I2 => sig00000287,
      I3 => sig000006d1,
      I4 => sig00000288,
      I5 => sig000006d1,
      O => sig0000028c
    );
  blk000001c6 : LUT6
    generic map(
      INIT => X"9009000000009009"
    )
    port map (
      I0 => sig00000283,
      I1 => sig000006d1,
      I2 => sig00000284,
      I3 => sig000008b6,
      I4 => sig00000285,
      I5 => sig000006d1,
      O => sig0000028d
    );
  blk000001c7 : MUXCY
    port map (
      CI => sig0000028f,
      DI => sig000008b6,
      S => sig0000028c,
      O => sig0000028e
    );
  blk000001c8 : MUXCY
    port map (
      CI => sig000006d1,
      DI => sig000008b6,
      S => sig0000028d,
      O => sig0000028f
    );
  blk000001c9 : XORCY
    port map (
      CI => sig0000028e,
      LI => sig000008b6,
      O => sig00000290
    );
  blk000001ca : MUXCY
    port map (
      CI => sig000006d1,
      DI => sig000008b6,
      S => sig00000298,
      O => sig00000299
    );
  blk000001cb : XORCY
    port map (
      CI => sig0000029b,
      LI => sig000008b6,
      O => sig0000029a
    );
  blk000001cc : MUXCY
    port map (
      CI => sig0000029c,
      DI => sig000008b6,
      S => sig0000029e,
      O => sig0000029b
    );
  blk000001cd : LUT3
    generic map(
      INIT => X"AE"
    )
    port map (
      I0 => sig00000112,
      I1 => sig0000029f,
      I2 => sig000002a0,
      O => sig0000029d
    );
  blk000001ce : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => sig0000029e,
      D => sig00000291,
      R => sig000008b6,
      Q => sig000002a0
    );
  blk000001cf : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => sig0000029e,
      D => sig00000290,
      R => sig000008b6,
      Q => sig00000291
    );
  blk000001d0 : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => sig0000029a,
      R => sig000008b6,
      Q => sig00000282
    );
  blk000001d1 : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => sig0000029d,
      R => sig000008b6,
      Q => sig0000029f
    );
  blk000001e9 : LUT6
    generic map(
      INIT => X"9009000000009009"
    )
    port map (
      I0 => sig0000027f,
      I1 => sig000008b6,
      I2 => sig00000280,
      I3 => sig000008b6,
      I4 => sig00000281,
      I5 => sig000008b6,
      O => sig000002a1
    );
  blk000001ea : LUT6
    generic map(
      INIT => X"9009000000009009"
    )
    port map (
      I0 => sig0000027c,
      I1 => sig000008b6,
      I2 => sig0000027d,
      I3 => sig000006d1,
      I4 => sig0000027e,
      I5 => sig000006d1,
      O => sig000002a2
    );
  blk000001eb : MUXCY
    port map (
      CI => sig000002a3,
      DI => sig000008b6,
      S => sig000002a1,
      O => sig000002b4
    );
  blk000001ec : MUXCY
    port map (
      CI => sig000006d1,
      DI => sig000008b6,
      S => sig000002a2,
      O => sig000002a3
    );
  blk000001ed : LUT6
    generic map(
      INIT => X"9009000000009009"
    )
    port map (
      I0 => sig0000027f,
      I1 => sig000006d1,
      I2 => sig00000280,
      I3 => sig000006d1,
      I4 => sig00000281,
      I5 => sig000006d1,
      O => sig000002a4
    );
  blk000001ee : LUT6
    generic map(
      INIT => X"9009000000009009"
    )
    port map (
      I0 => sig0000027c,
      I1 => sig000006d1,
      I2 => sig0000027d,
      I3 => sig000008b6,
      I4 => sig0000027e,
      I5 => sig000006d1,
      O => sig000002a5
    );
  blk000001ef : MUXCY
    port map (
      CI => sig000002a7,
      DI => sig000008b6,
      S => sig000002a4,
      O => sig000002a6
    );
  blk000001f0 : MUXCY
    port map (
      CI => sig000006d1,
      DI => sig000008b6,
      S => sig000002a5,
      O => sig000002a7
    );
  blk000001f1 : XORCY
    port map (
      CI => sig000002a6,
      LI => sig000008b6,
      O => sig000002a8
    );
  blk000001f2 : MUXCY
    port map (
      CI => sig000006d1,
      DI => sig000008b6,
      S => sig000002b0,
      O => sig000002b1
    );
  blk000001f3 : XORCY
    port map (
      CI => sig000002b3,
      LI => sig000008b6,
      O => sig000002b2
    );
  blk000001f4 : MUXCY
    port map (
      CI => sig000002b4,
      DI => sig000008b6,
      S => sig000002b6,
      O => sig000002b3
    );
  blk000001f5 : LUT3
    generic map(
      INIT => X"AE"
    )
    port map (
      I0 => sig00000282,
      I1 => sig000002b7,
      I2 => sig000002b8,
      O => sig000002b5
    );
  blk000001f6 : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => sig000002b6,
      D => sig000002a9,
      R => sig000008b6,
      Q => sig000002b8
    );
  blk000001f7 : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => sig000002b6,
      D => sig000002a8,
      R => sig000008b6,
      Q => sig000002a9
    );
  blk000001f8 : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => sig000002b2,
      R => sig000008b6,
      Q => sig0000027b
    );
  blk000001f9 : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => sig000002b5,
      R => sig000008b6,
      Q => sig000002b7
    );
  blk00000238 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => sig0000030c,
      Q => sig0000030b
    );
  blk00000239 : SRL16E
    generic map(
      INIT => X"0000"
    )
    port map (
      A0 => sig000006d1,
      A1 => sig000006d1,
      A2 => sig000008b6,
      A3 => sig000008b6,
      CE => ce,
      CLK => clk,
      D => sig00000136,
      Q => sig00000325
    );
  blk0000023a : SRL16E
    generic map(
      INIT => X"0000"
    )
    port map (
      A0 => sig000006d1,
      A1 => sig000006d1,
      A2 => sig000008b6,
      A3 => sig000008b6,
      CE => ce,
      CLK => clk,
      D => sig00000137,
      Q => sig00000326
    );
  blk0000023b : SRL16E
    generic map(
      INIT => X"0000"
    )
    port map (
      A0 => sig000006d1,
      A1 => sig000006d1,
      A2 => sig000008b6,
      A3 => sig000008b6,
      CE => ce,
      CLK => clk,
      D => sig00000138,
      Q => sig00000327
    );
  blk0000023c : SRL16E
    generic map(
      INIT => X"0000"
    )
    port map (
      A0 => sig000006d1,
      A1 => sig000006d1,
      A2 => sig000008b6,
      A3 => sig000008b6,
      CE => ce,
      CLK => clk,
      D => sig00000139,
      Q => sig00000328
    );
  blk0000023d : SRL16E
    generic map(
      INIT => X"0000"
    )
    port map (
      A0 => sig000006d1,
      A1 => sig000006d1,
      A2 => sig000008b6,
      A3 => sig000008b6,
      CE => ce,
      CLK => clk,
      D => sig0000013a,
      Q => sig00000329
    );
  blk0000023e : SRL16E
    generic map(
      INIT => X"0000"
    )
    port map (
      A0 => sig000006d1,
      A1 => sig000006d1,
      A2 => sig000008b6,
      A3 => sig000008b6,
      CE => ce,
      CLK => clk,
      D => sig0000013b,
      Q => sig0000032a
    );
  blk0000023f : SRL16E
    generic map(
      INIT => X"0000"
    )
    port map (
      A0 => sig000006d1,
      A1 => sig000006d1,
      A2 => sig000008b6,
      A3 => sig000008b6,
      CE => ce,
      CLK => clk,
      D => sig0000013c,
      Q => sig0000032b
    );
  blk00000240 : SRL16E
    generic map(
      INIT => X"0000"
    )
    port map (
      A0 => sig000006d1,
      A1 => sig000006d1,
      A2 => sig000008b6,
      A3 => sig000008b6,
      CE => ce,
      CLK => clk,
      D => sig0000013d,
      Q => sig0000032c
    );
  blk00000241 : SRL16E
    generic map(
      INIT => X"0000"
    )
    port map (
      A0 => sig000006d1,
      A1 => sig000006d1,
      A2 => sig000008b6,
      A3 => sig000008b6,
      CE => ce,
      CLK => clk,
      D => sig0000013e,
      Q => sig0000032d
    );
  blk00000242 : SRL16E
    generic map(
      INIT => X"0000"
    )
    port map (
      A0 => sig000006d1,
      A1 => sig000006d1,
      A2 => sig000008b6,
      A3 => sig000008b6,
      CE => ce,
      CLK => clk,
      D => sig0000013f,
      Q => sig0000032e
    );
  blk00000243 : SRL16E
    generic map(
      INIT => X"0000"
    )
    port map (
      A0 => sig000006d1,
      A1 => sig000006d1,
      A2 => sig000008b6,
      A3 => sig000008b6,
      CE => ce,
      CLK => clk,
      D => sig00000140,
      Q => sig0000032f
    );
  blk00000244 : SRL16E
    generic map(
      INIT => X"0000"
    )
    port map (
      A0 => sig000006d1,
      A1 => sig000006d1,
      A2 => sig000008b6,
      A3 => sig000008b6,
      CE => ce,
      CLK => clk,
      D => sig00000141,
      Q => sig00000330
    );
  blk00000245 : SRL16E
    generic map(
      INIT => X"0000"
    )
    port map (
      A0 => sig000006d1,
      A1 => sig000006d1,
      A2 => sig000008b6,
      A3 => sig000008b6,
      CE => ce,
      CLK => clk,
      D => sig00000141,
      Q => sig00000331
    );
  blk00000246 : MUXF7
    port map (
      I0 => sig00000325,
      I1 => sig00000ef7,
      S => sig0000030b,
      O => sig00000332
    );
  blk00000247 : MUXF7
    port map (
      I0 => sig00000326,
      I1 => sig00000ef8,
      S => sig0000030b,
      O => sig00000333
    );
  blk00000248 : MUXF7
    port map (
      I0 => sig00000327,
      I1 => sig00000ef9,
      S => sig0000030b,
      O => sig00000334
    );
  blk00000249 : MUXF7
    port map (
      I0 => sig00000328,
      I1 => sig00000efa,
      S => sig0000030b,
      O => sig00000335
    );
  blk0000024a : MUXF7
    port map (
      I0 => sig00000329,
      I1 => sig00000efb,
      S => sig0000030b,
      O => sig00000336
    );
  blk0000024b : MUXF7
    port map (
      I0 => sig0000032a,
      I1 => sig00000efc,
      S => sig0000030b,
      O => sig00000337
    );
  blk0000024c : MUXF7
    port map (
      I0 => sig0000032b,
      I1 => sig00000efd,
      S => sig0000030b,
      O => sig00000338
    );
  blk0000024d : MUXF7
    port map (
      I0 => sig0000032c,
      I1 => sig00000efe,
      S => sig0000030b,
      O => sig00000339
    );
  blk0000024e : MUXF7
    port map (
      I0 => sig0000032d,
      I1 => sig00000eff,
      S => sig0000030b,
      O => sig0000033a
    );
  blk0000024f : MUXF7
    port map (
      I0 => sig0000032e,
      I1 => sig00000f00,
      S => sig0000030b,
      O => sig0000033b
    );
  blk00000250 : MUXF7
    port map (
      I0 => sig0000032f,
      I1 => sig00000f01,
      S => sig0000030b,
      O => sig0000033c
    );
  blk00000251 : MUXF7
    port map (
      I0 => sig00000330,
      I1 => sig00000f02,
      S => sig0000030b,
      O => sig0000033d
    );
  blk00000252 : MUXF7
    port map (
      I0 => sig00000331,
      I1 => sig00000f03,
      S => sig0000030b,
      O => sig0000033e
    );
  blk00000253 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => sig00000332,
      Q => sig000002fe
    );
  blk00000254 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => sig00000333,
      Q => sig000002ff
    );
  blk00000255 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => sig00000334,
      Q => sig00000300
    );
  blk00000256 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => sig00000335,
      Q => sig00000301
    );
  blk00000257 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => sig00000336,
      Q => sig00000302
    );
  blk00000258 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => sig00000337,
      Q => sig00000303
    );
  blk00000259 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => sig00000338,
      Q => sig00000304
    );
  blk0000025a : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => sig00000339,
      Q => sig00000305
    );
  blk0000025b : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => sig0000033a,
      Q => sig00000306
    );
  blk0000025c : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => sig0000033b,
      Q => sig00000307
    );
  blk0000025d : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => sig0000033c,
      Q => sig00000308
    );
  blk0000025e : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => sig0000033d,
      Q => sig00000309
    );
  blk0000025f : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => sig0000033e,
      Q => sig0000030a
    );
  blk00000260 : SRL16E
    generic map(
      INIT => X"0000"
    )
    port map (
      A0 => sig000006d1,
      A1 => sig000006d1,
      A2 => sig000008b6,
      A3 => sig000008b6,
      CE => ce,
      CLK => clk,
      D => sig0000012a,
      Q => sig0000033f
    );
  blk00000261 : SRL16E
    generic map(
      INIT => X"0000"
    )
    port map (
      A0 => sig000006d1,
      A1 => sig000006d1,
      A2 => sig000008b6,
      A3 => sig000008b6,
      CE => ce,
      CLK => clk,
      D => sig0000012b,
      Q => sig00000340
    );
  blk00000262 : SRL16E
    generic map(
      INIT => X"0000"
    )
    port map (
      A0 => sig000006d1,
      A1 => sig000006d1,
      A2 => sig000008b6,
      A3 => sig000008b6,
      CE => ce,
      CLK => clk,
      D => sig0000012c,
      Q => sig00000341
    );
  blk00000263 : SRL16E
    generic map(
      INIT => X"0000"
    )
    port map (
      A0 => sig000006d1,
      A1 => sig000006d1,
      A2 => sig000008b6,
      A3 => sig000008b6,
      CE => ce,
      CLK => clk,
      D => sig0000012d,
      Q => sig00000342
    );
  blk00000264 : SRL16E
    generic map(
      INIT => X"0000"
    )
    port map (
      A0 => sig000006d1,
      A1 => sig000006d1,
      A2 => sig000008b6,
      A3 => sig000008b6,
      CE => ce,
      CLK => clk,
      D => sig0000012e,
      Q => sig00000343
    );
  blk00000265 : SRL16E
    generic map(
      INIT => X"0000"
    )
    port map (
      A0 => sig000006d1,
      A1 => sig000006d1,
      A2 => sig000008b6,
      A3 => sig000008b6,
      CE => ce,
      CLK => clk,
      D => sig0000012f,
      Q => sig00000344
    );
  blk00000266 : SRL16E
    generic map(
      INIT => X"0000"
    )
    port map (
      A0 => sig000006d1,
      A1 => sig000006d1,
      A2 => sig000008b6,
      A3 => sig000008b6,
      CE => ce,
      CLK => clk,
      D => sig00000130,
      Q => sig00000345
    );
  blk00000267 : SRL16E
    generic map(
      INIT => X"0000"
    )
    port map (
      A0 => sig000006d1,
      A1 => sig000006d1,
      A2 => sig000008b6,
      A3 => sig000008b6,
      CE => ce,
      CLK => clk,
      D => sig00000131,
      Q => sig00000346
    );
  blk00000268 : SRL16E
    generic map(
      INIT => X"0000"
    )
    port map (
      A0 => sig000006d1,
      A1 => sig000006d1,
      A2 => sig000008b6,
      A3 => sig000008b6,
      CE => ce,
      CLK => clk,
      D => sig00000132,
      Q => sig00000347
    );
  blk00000269 : SRL16E
    generic map(
      INIT => X"0000"
    )
    port map (
      A0 => sig000006d1,
      A1 => sig000006d1,
      A2 => sig000008b6,
      A3 => sig000008b6,
      CE => ce,
      CLK => clk,
      D => sig00000133,
      Q => sig00000348
    );
  blk0000026a : SRL16E
    generic map(
      INIT => X"0000"
    )
    port map (
      A0 => sig000006d1,
      A1 => sig000006d1,
      A2 => sig000008b6,
      A3 => sig000008b6,
      CE => ce,
      CLK => clk,
      D => sig00000134,
      Q => sig00000349
    );
  blk0000026b : SRL16E
    generic map(
      INIT => X"0000"
    )
    port map (
      A0 => sig000006d1,
      A1 => sig000006d1,
      A2 => sig000008b6,
      A3 => sig000008b6,
      CE => ce,
      CLK => clk,
      D => sig00000135,
      Q => sig0000034a
    );
  blk0000026c : SRL16E
    generic map(
      INIT => X"0000"
    )
    port map (
      A0 => sig000006d1,
      A1 => sig000006d1,
      A2 => sig000008b6,
      A3 => sig000008b6,
      CE => ce,
      CLK => clk,
      D => sig00000135,
      Q => sig0000034b
    );
  blk0000026d : MUXF7
    port map (
      I0 => sig0000033f,
      I1 => sig00000f04,
      S => sig0000030b,
      O => sig0000034c
    );
  blk0000026e : MUXF7
    port map (
      I0 => sig00000340,
      I1 => sig00000f05,
      S => sig0000030b,
      O => sig0000034d
    );
  blk0000026f : MUXF7
    port map (
      I0 => sig00000341,
      I1 => sig00000f06,
      S => sig0000030b,
      O => sig0000034e
    );
  blk00000270 : MUXF7
    port map (
      I0 => sig00000342,
      I1 => sig00000f07,
      S => sig0000030b,
      O => sig0000034f
    );
  blk00000271 : MUXF7
    port map (
      I0 => sig00000343,
      I1 => sig00000f08,
      S => sig0000030b,
      O => sig00000350
    );
  blk00000272 : MUXF7
    port map (
      I0 => sig00000344,
      I1 => sig00000f09,
      S => sig0000030b,
      O => sig00000351
    );
  blk00000273 : MUXF7
    port map (
      I0 => sig00000345,
      I1 => sig00000f0a,
      S => sig0000030b,
      O => sig00000352
    );
  blk00000274 : MUXF7
    port map (
      I0 => sig00000346,
      I1 => sig00000f0b,
      S => sig0000030b,
      O => sig00000353
    );
  blk00000275 : MUXF7
    port map (
      I0 => sig00000347,
      I1 => sig00000f0c,
      S => sig0000030b,
      O => sig00000354
    );
  blk00000276 : MUXF7
    port map (
      I0 => sig00000348,
      I1 => sig00000f0d,
      S => sig0000030b,
      O => sig00000355
    );
  blk00000277 : MUXF7
    port map (
      I0 => sig00000349,
      I1 => sig00000f0e,
      S => sig0000030b,
      O => sig00000356
    );
  blk00000278 : MUXF7
    port map (
      I0 => sig0000034a,
      I1 => sig00000f0f,
      S => sig0000030b,
      O => sig00000357
    );
  blk00000279 : MUXF7
    port map (
      I0 => sig0000034b,
      I1 => sig00000f10,
      S => sig0000030b,
      O => sig00000358
    );
  blk0000027a : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => sig0000034c,
      Q => sig000002f1
    );
  blk0000027b : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => sig0000034d,
      Q => sig000002f2
    );
  blk0000027c : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => sig0000034e,
      Q => sig000002f3
    );
  blk0000027d : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => sig0000034f,
      Q => sig000002f4
    );
  blk0000027e : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => sig00000350,
      Q => sig000002f5
    );
  blk0000027f : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => sig00000351,
      Q => sig000002f6
    );
  blk00000280 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => sig00000352,
      Q => sig000002f7
    );
  blk00000281 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => sig00000353,
      Q => sig000002f8
    );
  blk00000282 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => sig00000354,
      Q => sig000002f9
    );
  blk00000283 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => sig00000355,
      Q => sig000002fa
    );
  blk00000284 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => sig00000356,
      Q => sig000002fb
    );
  blk00000285 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => sig00000357,
      Q => sig000002fc
    );
  blk00000286 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => sig00000358,
      Q => sig000002fd
    );
  blk000003f3 : MUXCY
    port map (
      CI => sig000003ba,
      DI => sig000008b6,
      S => sig00000391,
      O => sig0000039f
    );
  blk000003f4 : XORCY
    port map (
      CI => sig000003ba,
      LI => sig00000391,
      O => sig000003a0
    );
  blk000003f5 : MUXCY
    port map (
      CI => sig0000039f,
      DI => sig000008b6,
      S => sig00000392,
      O => sig000003a1
    );
  blk000003f6 : XORCY
    port map (
      CI => sig0000039f,
      LI => sig00000392,
      O => sig000003a2
    );
  blk000003f7 : MUXCY
    port map (
      CI => sig000003a1,
      DI => sig000008b6,
      S => sig00000393,
      O => sig000003a3
    );
  blk000003f8 : XORCY
    port map (
      CI => sig000003a1,
      LI => sig00000393,
      O => sig000003a4
    );
  blk000003f9 : MUXCY
    port map (
      CI => sig000003a3,
      DI => sig000008b6,
      S => sig00000394,
      O => sig000003a5
    );
  blk000003fa : XORCY
    port map (
      CI => sig000003a3,
      LI => sig00000394,
      O => sig000003a6
    );
  blk000003fb : MUXCY
    port map (
      CI => sig000003a5,
      DI => sig000008b6,
      S => sig00000395,
      O => sig000003a7
    );
  blk000003fc : XORCY
    port map (
      CI => sig000003a5,
      LI => sig00000395,
      O => sig000003a8
    );
  blk000003fd : MUXCY
    port map (
      CI => sig000003a7,
      DI => sig000008b6,
      S => sig00000396,
      O => sig000003a9
    );
  blk000003fe : XORCY
    port map (
      CI => sig000003a7,
      LI => sig00000396,
      O => sig000003aa
    );
  blk000003ff : MUXCY
    port map (
      CI => sig000003a9,
      DI => sig000008b6,
      S => sig00000397,
      O => sig000003ab
    );
  blk00000400 : XORCY
    port map (
      CI => sig000003a9,
      LI => sig00000397,
      O => sig000003ac
    );
  blk00000401 : MUXCY
    port map (
      CI => sig000003ab,
      DI => sig000008b6,
      S => sig00000398,
      O => sig000003ad
    );
  blk00000402 : XORCY
    port map (
      CI => sig000003ab,
      LI => sig00000398,
      O => sig000003ae
    );
  blk00000403 : MUXCY
    port map (
      CI => sig000003ad,
      DI => sig000008b6,
      S => sig00000399,
      O => sig000003af
    );
  blk00000404 : XORCY
    port map (
      CI => sig000003ad,
      LI => sig00000399,
      O => sig000003b0
    );
  blk00000405 : MUXCY
    port map (
      CI => sig000003af,
      DI => sig000008b6,
      S => sig0000039a,
      O => sig000003b1
    );
  blk00000406 : XORCY
    port map (
      CI => sig000003af,
      LI => sig0000039a,
      O => sig000003b2
    );
  blk00000407 : MUXCY
    port map (
      CI => sig000003b1,
      DI => sig000008b6,
      S => sig0000039b,
      O => sig000003b3
    );
  blk00000408 : XORCY
    port map (
      CI => sig000003b1,
      LI => sig0000039b,
      O => sig000003b4
    );
  blk00000409 : MUXCY
    port map (
      CI => sig000003b3,
      DI => sig000008b6,
      S => sig0000039c,
      O => sig000003b5
    );
  blk0000040a : XORCY
    port map (
      CI => sig000003b3,
      LI => sig0000039c,
      O => sig000003b6
    );
  blk0000040b : MUXCY
    port map (
      CI => sig000003b5,
      DI => sig000008b6,
      S => sig00000eee,
      O => sig000003b7
    );
  blk0000040c : XORCY
    port map (
      CI => sig000003b5,
      LI => sig00000eee,
      O => sig000003b8
    );
  blk0000040d : MUXCY
    port map (
      CI => sig000003b7,
      DI => sig000008b6,
      S => sig0000039d,
      O => NLW_blk0000040d_O_UNCONNECTED
    );
  blk0000040e : XORCY
    port map (
      CI => sig000003b7,
      LI => sig0000039d,
      O => sig000003b9
    );
  blk0000040f : MUXCY
    port map (
      CI => sig000006d1,
      DI => sig000008b6,
      S => sig0000039e,
      O => sig000003ba
    );
  blk00000410 : MUXCY
    port map (
      CI => sig000003e4,
      DI => sig000008b6,
      S => sig000003bb,
      O => sig000003c9
    );
  blk00000411 : XORCY
    port map (
      CI => sig000003e4,
      LI => sig000003bb,
      O => sig000003ca
    );
  blk00000412 : MUXCY
    port map (
      CI => sig000003c9,
      DI => sig000008b6,
      S => sig000003bc,
      O => sig000003cb
    );
  blk00000413 : XORCY
    port map (
      CI => sig000003c9,
      LI => sig000003bc,
      O => sig000003cc
    );
  blk00000414 : MUXCY
    port map (
      CI => sig000003cb,
      DI => sig000008b6,
      S => sig000003bd,
      O => sig000003cd
    );
  blk00000415 : XORCY
    port map (
      CI => sig000003cb,
      LI => sig000003bd,
      O => sig000003ce
    );
  blk00000416 : MUXCY
    port map (
      CI => sig000003cd,
      DI => sig000008b6,
      S => sig000003be,
      O => sig000003cf
    );
  blk00000417 : XORCY
    port map (
      CI => sig000003cd,
      LI => sig000003be,
      O => sig000003d0
    );
  blk00000418 : MUXCY
    port map (
      CI => sig000003cf,
      DI => sig000008b6,
      S => sig000003bf,
      O => sig000003d1
    );
  blk00000419 : XORCY
    port map (
      CI => sig000003cf,
      LI => sig000003bf,
      O => sig000003d2
    );
  blk0000041a : MUXCY
    port map (
      CI => sig000003d1,
      DI => sig000008b6,
      S => sig000003c0,
      O => sig000003d3
    );
  blk0000041b : XORCY
    port map (
      CI => sig000003d1,
      LI => sig000003c0,
      O => sig000003d4
    );
  blk0000041c : MUXCY
    port map (
      CI => sig000003d3,
      DI => sig000008b6,
      S => sig000003c1,
      O => sig000003d5
    );
  blk0000041d : XORCY
    port map (
      CI => sig000003d3,
      LI => sig000003c1,
      O => sig000003d6
    );
  blk0000041e : MUXCY
    port map (
      CI => sig000003d5,
      DI => sig000008b6,
      S => sig000003c2,
      O => sig000003d7
    );
  blk0000041f : XORCY
    port map (
      CI => sig000003d5,
      LI => sig000003c2,
      O => sig000003d8
    );
  blk00000420 : MUXCY
    port map (
      CI => sig000003d7,
      DI => sig000008b6,
      S => sig000003c3,
      O => sig000003d9
    );
  blk00000421 : XORCY
    port map (
      CI => sig000003d7,
      LI => sig000003c3,
      O => sig000003da
    );
  blk00000422 : MUXCY
    port map (
      CI => sig000003d9,
      DI => sig000008b6,
      S => sig000003c4,
      O => sig000003db
    );
  blk00000423 : XORCY
    port map (
      CI => sig000003d9,
      LI => sig000003c4,
      O => sig000003dc
    );
  blk00000424 : MUXCY
    port map (
      CI => sig000003db,
      DI => sig000008b6,
      S => sig000003c5,
      O => sig000003dd
    );
  blk00000425 : XORCY
    port map (
      CI => sig000003db,
      LI => sig000003c5,
      O => sig000003de
    );
  blk00000426 : MUXCY
    port map (
      CI => sig000003dd,
      DI => sig000008b6,
      S => sig000003c6,
      O => sig000003df
    );
  blk00000427 : XORCY
    port map (
      CI => sig000003dd,
      LI => sig000003c6,
      O => sig000003e0
    );
  blk00000428 : MUXCY
    port map (
      CI => sig000003df,
      DI => sig000008b6,
      S => sig00000eef,
      O => sig000003e1
    );
  blk00000429 : XORCY
    port map (
      CI => sig000003df,
      LI => sig00000eef,
      O => sig000003e2
    );
  blk0000042a : MUXCY
    port map (
      CI => sig000003e1,
      DI => sig000008b6,
      S => sig000003c7,
      O => NLW_blk0000042a_O_UNCONNECTED
    );
  blk0000042b : XORCY
    port map (
      CI => sig000003e1,
      LI => sig000003c7,
      O => sig000003e3
    );
  blk0000042c : MUXCY
    port map (
      CI => sig000006d1,
      DI => sig000008b6,
      S => sig000003c8,
      O => sig000003e4
    );
  blk0000042d : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => sig00000366,
      R => sig000008b6,
      Q => sig00000448
    );
  blk0000042e : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => sig00000365,
      R => sig000008b6,
      Q => sig00000449
    );
  blk0000042f : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => sig00000364,
      R => sig000008b6,
      Q => sig0000044a
    );
  blk00000430 : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => sig00000363,
      R => sig000008b6,
      Q => sig0000044b
    );
  blk00000431 : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => sig00000362,
      R => sig000008b6,
      Q => sig0000044c
    );
  blk00000432 : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => sig00000361,
      R => sig000008b6,
      Q => sig0000044d
    );
  blk00000433 : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => sig00000360,
      R => sig000008b6,
      Q => sig0000044e
    );
  blk00000434 : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => sig0000035f,
      R => sig000008b6,
      Q => sig0000044f
    );
  blk00000435 : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => sig0000035e,
      R => sig000008b6,
      Q => sig00000450
    );
  blk00000436 : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => sig0000035d,
      R => sig000008b6,
      Q => sig00000451
    );
  blk00000437 : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => sig0000035c,
      R => sig000008b6,
      Q => sig00000452
    );
  blk00000438 : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => sig0000035b,
      R => sig000008b6,
      Q => sig00000453
    );
  blk00000439 : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => sig0000035a,
      R => sig000008b6,
      Q => sig00000454
    );
  blk0000043a : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => sig00000359,
      R => sig000008b6,
      Q => sig00000455
    );
  blk0000043b : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => sig00000374,
      R => sig000008b6,
      Q => sig0000043a
    );
  blk0000043c : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => sig00000373,
      R => sig000008b6,
      Q => sig0000043b
    );
  blk0000043d : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => sig00000372,
      R => sig000008b6,
      Q => sig0000043c
    );
  blk0000043e : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => sig00000371,
      R => sig000008b6,
      Q => sig0000043d
    );
  blk0000043f : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => sig00000370,
      R => sig000008b6,
      Q => sig0000043e
    );
  blk00000440 : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => sig0000036f,
      R => sig000008b6,
      Q => sig0000043f
    );
  blk00000441 : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => sig0000036e,
      R => sig000008b6,
      Q => sig00000440
    );
  blk00000442 : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => sig0000036d,
      R => sig000008b6,
      Q => sig00000441
    );
  blk00000443 : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => sig0000036c,
      R => sig000008b6,
      Q => sig00000442
    );
  blk00000444 : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => sig0000036b,
      R => sig000008b6,
      Q => sig00000443
    );
  blk00000445 : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => sig0000036a,
      R => sig000008b6,
      Q => sig00000444
    );
  blk00000446 : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => sig00000369,
      R => sig000008b6,
      Q => sig00000445
    );
  blk00000447 : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => sig00000368,
      R => sig000008b6,
      Q => sig00000446
    );
  blk00000448 : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => sig00000367,
      R => sig000008b6,
      Q => sig00000447
    );
  blk00000449 : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => sig00000382,
      R => sig000008b6,
      Q => sig00000402
    );
  blk0000044a : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => sig00000381,
      R => sig000008b6,
      Q => sig00000403
    );
  blk0000044b : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => sig00000380,
      R => sig000008b6,
      Q => sig00000404
    );
  blk0000044c : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => sig0000037f,
      R => sig000008b6,
      Q => sig00000405
    );
  blk0000044d : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => sig0000037e,
      R => sig000008b6,
      Q => sig00000406
    );
  blk0000044e : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => sig0000037d,
      R => sig000008b6,
      Q => sig00000407
    );
  blk0000044f : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => sig0000037c,
      R => sig000008b6,
      Q => sig00000408
    );
  blk00000450 : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => sig0000037b,
      R => sig000008b6,
      Q => sig00000409
    );
  blk00000451 : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => sig0000037a,
      R => sig000008b6,
      Q => sig0000040a
    );
  blk00000452 : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => sig00000379,
      R => sig000008b6,
      Q => sig0000040b
    );
  blk00000453 : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => sig00000378,
      R => sig000008b6,
      Q => sig0000040c
    );
  blk00000454 : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => sig00000377,
      R => sig000008b6,
      Q => sig0000040d
    );
  blk00000455 : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => sig00000376,
      R => sig000008b6,
      Q => sig0000040e
    );
  blk00000456 : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => sig00000375,
      R => sig000008b6,
      Q => sig0000040f
    );
  blk00000457 : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => sig00000390,
      R => sig000008b6,
      Q => sig00000233
    );
  blk00000458 : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => sig0000038f,
      R => sig000008b6,
      Q => sig00000234
    );
  blk00000459 : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => sig0000038e,
      R => sig000008b6,
      Q => sig00000235
    );
  blk0000045a : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => sig0000038d,
      R => sig000008b6,
      Q => sig00000236
    );
  blk0000045b : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => sig0000038c,
      R => sig000008b6,
      Q => sig00000237
    );
  blk0000045c : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => sig0000038b,
      R => sig000008b6,
      Q => sig00000238
    );
  blk0000045d : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => sig0000038a,
      R => sig000008b6,
      Q => sig00000239
    );
  blk0000045e : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => sig00000389,
      R => sig000008b6,
      Q => sig0000023a
    );
  blk0000045f : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => sig00000388,
      R => sig000008b6,
      Q => sig0000023b
    );
  blk00000460 : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => sig00000387,
      R => sig000008b6,
      Q => sig0000023c
    );
  blk00000461 : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => sig00000386,
      R => sig000008b6,
      Q => sig0000023d
    );
  blk00000462 : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => sig00000385,
      R => sig000008b6,
      Q => sig0000023e
    );
  blk00000463 : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => sig00000384,
      R => sig000008b6,
      Q => sig0000023f
    );
  blk00000464 : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => sig00000383,
      R => sig000008b6,
      Q => sig00000240
    );
  blk00000465 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => sig000003a0,
      Q => sig00000472
    );
  blk00000466 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => sig000003a2,
      Q => sig00000473
    );
  blk00000467 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => sig000003a4,
      Q => sig00000474
    );
  blk00000468 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => sig000003a6,
      Q => sig00000475
    );
  blk00000469 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => sig000003a8,
      Q => sig00000476
    );
  blk0000046a : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => sig000003aa,
      Q => sig00000477
    );
  blk0000046b : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => sig000003ac,
      Q => sig00000478
    );
  blk0000046c : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => sig000003ae,
      Q => sig00000479
    );
  blk0000046d : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => sig000003b0,
      Q => sig0000047a
    );
  blk0000046e : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => sig000003b2,
      Q => sig0000047b
    );
  blk0000046f : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => sig000003b4,
      Q => sig0000047c
    );
  blk00000470 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => sig000003b6,
      Q => sig0000047d
    );
  blk00000471 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => sig000003b8,
      Q => sig0000047e
    );
  blk00000472 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => sig000003b9,
      Q => sig0000047f
    );
  blk00000473 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => sig000003ca,
      Q => sig00000480
    );
  blk00000474 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => sig000003cc,
      Q => sig00000481
    );
  blk00000475 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => sig000003ce,
      Q => sig00000482
    );
  blk00000476 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => sig000003d0,
      Q => sig00000483
    );
  blk00000477 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => sig000003d2,
      Q => sig00000484
    );
  blk00000478 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => sig000003d4,
      Q => sig00000485
    );
  blk00000479 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => sig000003d6,
      Q => sig00000486
    );
  blk0000047a : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => sig000003d8,
      Q => sig00000487
    );
  blk0000047b : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => sig000003da,
      Q => sig00000488
    );
  blk0000047c : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => sig000003dc,
      Q => sig00000489
    );
  blk0000047d : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => sig000003de,
      Q => sig0000048a
    );
  blk0000047e : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => sig000003e0,
      Q => sig0000048b
    );
  blk0000047f : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => sig000003e2,
      Q => sig0000048c
    );
  blk00000480 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => sig000003e3,
      Q => sig0000048d
    );
  blk00000481 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => sig00000259,
      Q => sig00000493
    );
  blk00000482 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => sig000003e5,
      Q => sig0000048e
    );
  blk00000483 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => sig0000024f,
      Q => sig00000492
    );
  blk00000484 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => sig0000048d,
      Q => sig000003f3
    );
  blk00000485 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => sig0000048c,
      Q => sig000003f2
    );
  blk00000486 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => sig0000048b,
      Q => sig000003f1
    );
  blk00000487 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => sig0000048a,
      Q => sig000003f0
    );
  blk00000488 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => sig00000489,
      Q => sig000003ef
    );
  blk00000489 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => sig00000488,
      Q => sig000003ee
    );
  blk0000048a : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => sig00000487,
      Q => sig000003ed
    );
  blk0000048b : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => sig00000486,
      Q => sig000003ec
    );
  blk0000048c : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => sig00000485,
      Q => sig000003eb
    );
  blk0000048d : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => sig00000484,
      Q => sig000003ea
    );
  blk0000048e : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => sig00000483,
      Q => sig000003e9
    );
  blk0000048f : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => sig00000482,
      Q => sig000003e8
    );
  blk00000490 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => sig00000481,
      Q => sig000003e7
    );
  blk00000491 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => sig00000480,
      Q => sig000003e6
    );
  blk00000492 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => sig0000047f,
      Q => sig00000401
    );
  blk00000493 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => sig0000047e,
      Q => sig00000400
    );
  blk00000494 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => sig0000047d,
      Q => sig000003ff
    );
  blk00000495 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => sig0000047c,
      Q => sig000003fe
    );
  blk00000496 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => sig0000047b,
      Q => sig000003fd
    );
  blk00000497 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => sig0000047a,
      Q => sig000003fc
    );
  blk00000498 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => sig00000479,
      Q => sig000003fb
    );
  blk00000499 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => sig00000478,
      Q => sig000003fa
    );
  blk0000049a : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => sig00000477,
      Q => sig000003f9
    );
  blk0000049b : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => sig00000476,
      Q => sig000003f8
    );
  blk0000049c : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => sig00000475,
      Q => sig000003f7
    );
  blk0000049d : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => sig00000474,
      Q => sig000003f6
    );
  blk0000049e : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => sig00000473,
      Q => sig000003f5
    );
  blk0000049f : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => sig00000472,
      Q => sig000003f4
    );
  blk000005c7 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => sig0000022e,
      Q => sig000004a5
    );
  blk000005c8 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => sig0000022d,
      Q => sig000004a4
    );
  blk000005c9 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => sig00000232,
      Q => sig000004a9
    );
  blk000005ca : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => sig00000231,
      Q => sig000004a8
    );
  blk000005cb : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => sig00000230,
      Q => sig000004a7
    );
  blk000005cc : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => sig0000022f,
      Q => sig000004a6
    );
  blk000005e5 : LUT6
    generic map(
      INIT => X"FF00F0F0CCCCAAAA"
    )
    port map (
      I0 => sig000008b6,
      I1 => sig000008b6,
      I2 => sig000004a6,
      I3 => sig0000049e,
      I4 => sig000004a4,
      I5 => sig000004a5,
      O => sig000004aa
    );
  blk000005e6 : LUT6
    generic map(
      INIT => X"FF00F0F0CCCCAAAA"
    )
    port map (
      I0 => sig000008b6,
      I1 => sig000004a6,
      I2 => sig000004a7,
      I3 => sig0000049f,
      I4 => sig000004a4,
      I5 => sig000004a5,
      O => sig000004ab
    );
  blk000005e7 : LUT6
    generic map(
      INIT => X"FF00F0F0CCCCAAAA"
    )
    port map (
      I0 => sig000008b6,
      I1 => sig000004a7,
      I2 => sig000004a8,
      I3 => sig000004a0,
      I4 => sig000004a4,
      I5 => sig000004a5,
      O => sig000004ac
    );
  blk000005e8 : LUT6
    generic map(
      INIT => X"FF00F0F0CCCCAAAA"
    )
    port map (
      I0 => sig000008b6,
      I1 => sig000004a8,
      I2 => sig000004a9,
      I3 => sig000004a1,
      I4 => sig000004a4,
      I5 => sig000004a5,
      O => sig000004ad
    );
  blk000005e9 : LUT6
    generic map(
      INIT => X"FF00F0F0CCCCAAAA"
    )
    port map (
      I0 => sig000008b6,
      I1 => sig000004a9,
      I2 => sig000008b6,
      I3 => sig000004a2,
      I4 => sig000004a4,
      I5 => sig000004a5,
      O => sig000004ae
    );
  blk000005ea : LUT6
    generic map(
      INIT => X"FF00F0F0CCCCAAAA"
    )
    port map (
      I0 => sig000008b6,
      I1 => sig000008b6,
      I2 => sig000008b6,
      I3 => sig000004a3,
      I4 => sig000004a4,
      I5 => sig000004a5,
      O => sig000004af
    );
  blk000005eb : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => sig000004aa,
      R => sig000008b6,
      Q => sig00000499
    );
  blk000005ec : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => sig000004ab,
      R => sig000008b6,
      Q => sig0000049a
    );
  blk000005ed : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => sig000004ac,
      R => sig000008b6,
      Q => sig0000049b
    );
  blk000005ee : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => sig000004ad,
      R => sig000008b6,
      Q => sig0000049c
    );
  blk000005ef : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => sig000004ae,
      R => sig000008b6,
      Q => sig0000049d
    );
  blk000005f0 : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => sig000004af,
      R => sig000008b6,
      Q => sig00000498
    );
  blk00000655 : DSP48E
    generic map(
      ACASCREG => 2,
      ALUMODEREG => 0,
      AREG => 2,
      AUTORESET_PATTERN_DETECT => FALSE,
      AUTORESET_PATTERN_DETECT_OPTINV => "MATCH",
      A_INPUT => "DIRECT",
      BCASCREG => 2,
      BREG => 2,
      B_INPUT => "DIRECT",
      CARRYINREG => 0,
      CARRYINSELREG => 0,
      CREG => 1,
      MASK => X"000000000000",
      MREG => 1,
      MULTCARRYINREG => 0,
      OPMODEREG => 0,
      PATTERN => X"000000000000",
      PREG => 1,
      SEL_MASK => "MASK",
      SEL_PATTERN => "PATTERN",
      SEL_ROUNDING_MASK => "SEL_MASK",
      SIM_MODE => "SAFE",
      USE_MULT => "MULT_S",
      USE_PATTERN_DETECT => "NO_PATDET",
      USE_SIMD => "ONE48"
    )
    port map (
      CARRYIN => sig000008b6,
      CEA1 => ce,
      CEA2 => ce,
      CEB1 => ce,
      CEB2 => ce,
      CEC => ce,
      CECTRL => sig000008b6,
      CEP => ce,
      CEM => ce,
      CECARRYIN => sig000008b6,
      CEMULTCARRYIN => sig000008b6,
      CLK => clk,
      RSTA => sig000008b6,
      RSTB => sig000008b6,
      RSTC => sig000008b6,
      RSTCTRL => sig000008b6,
      RSTP => sig000008b6,
      RSTM => sig000008b6,
      RSTALLCARRYIN => sig000008b6,
      CEALUMODE => sig000008b6,
      RSTALUMODE => sig000008b6,
      PATTERNBDETECT => NLW_blk00000655_PATTERNBDETECT_UNCONNECTED,
      PATTERNDETECT => NLW_blk00000655_PATTERNDETECT_UNCONNECTED,
      OVERFLOW => NLW_blk00000655_OVERFLOW_UNCONNECTED,
      UNDERFLOW => NLW_blk00000655_UNDERFLOW_UNCONNECTED,
      CARRYCASCIN => sig000008b6,
      CARRYCASCOUT => NLW_blk00000655_CARRYCASCOUT_UNCONNECTED,
      MULTSIGNIN => sig000008b6,
      MULTSIGNOUT => NLW_blk00000655_MULTSIGNOUT_UNCONNECTED,
      A(29) => sig000008b6,
      A(28) => sig000008b6,
      A(27) => sig000008b6,
      A(26) => sig000008b6,
      A(25) => sig000008b6,
      A(24) => sig00000530,
      A(23) => sig00000530,
      A(22) => sig00000530,
      A(21) => sig00000530,
      A(20) => sig00000530,
      A(19) => sig00000530,
      A(18) => sig00000530,
      A(17) => sig00000530,
      A(16) => sig00000530,
      A(15) => sig00000530,
      A(14) => sig00000530,
      A(13) => sig00000530,
      A(12) => sig00000530,
      A(11) => sig0000053d,
      A(10) => sig0000053e,
      A(9) => sig0000053f,
      A(8) => sig00000540,
      A(7) => sig00000541,
      A(6) => sig00000542,
      A(5) => sig00000543,
      A(4) => sig00000544,
      A(3) => sig00000545,
      A(2) => sig00000546,
      A(1) => sig00000547,
      A(0) => sig00000548,
      PCIN(47) => sig000008b6,
      PCIN(46) => sig000008b6,
      PCIN(45) => sig000008b6,
      PCIN(44) => sig000008b6,
      PCIN(43) => sig000008b6,
      PCIN(42) => sig000008b6,
      PCIN(41) => sig000008b6,
      PCIN(40) => sig000008b6,
      PCIN(39) => sig000008b6,
      PCIN(38) => sig000008b6,
      PCIN(37) => sig000008b6,
      PCIN(36) => sig000008b6,
      PCIN(35) => sig000008b6,
      PCIN(34) => sig000008b6,
      PCIN(33) => sig000008b6,
      PCIN(32) => sig000008b6,
      PCIN(31) => sig000008b6,
      PCIN(30) => sig000008b6,
      PCIN(29) => sig000008b6,
      PCIN(28) => sig000008b6,
      PCIN(27) => sig000008b6,
      PCIN(26) => sig000008b6,
      PCIN(25) => sig000008b6,
      PCIN(24) => sig000008b6,
      PCIN(23) => sig000008b6,
      PCIN(22) => sig000008b6,
      PCIN(21) => sig000008b6,
      PCIN(20) => sig000008b6,
      PCIN(19) => sig000008b6,
      PCIN(18) => sig000008b6,
      PCIN(17) => sig000008b6,
      PCIN(16) => sig000008b6,
      PCIN(15) => sig000008b6,
      PCIN(14) => sig000008b6,
      PCIN(13) => sig000008b6,
      PCIN(12) => sig000008b6,
      PCIN(11) => sig000008b6,
      PCIN(10) => sig000008b6,
      PCIN(9) => sig000008b6,
      PCIN(8) => sig000008b6,
      PCIN(7) => sig000008b6,
      PCIN(6) => sig000008b6,
      PCIN(5) => sig000008b6,
      PCIN(4) => sig000008b6,
      PCIN(3) => sig000008b6,
      PCIN(2) => sig000008b6,
      PCIN(1) => sig000008b6,
      PCIN(0) => sig000008b6,
      B(17) => sig00000549,
      B(16) => sig00000549,
      B(15) => sig00000549,
      B(14) => sig00000549,
      B(13) => sig0000054d,
      B(12) => sig0000054e,
      B(11) => sig0000054f,
      B(10) => sig00000550,
      B(9) => sig00000551,
      B(8) => sig00000552,
      B(7) => sig00000553,
      B(6) => sig00000554,
      B(5) => sig00000555,
      B(4) => sig00000556,
      B(3) => sig00000557,
      B(2) => sig00000558,
      B(1) => sig00000559,
      B(0) => sig0000055a,
      C(47) => sig0000056a,
      C(46) => sig0000056a,
      C(45) => sig0000056a,
      C(44) => sig0000056a,
      C(43) => sig0000056a,
      C(42) => sig0000056a,
      C(41) => sig0000056a,
      C(40) => sig0000056a,
      C(39) => sig0000056a,
      C(38) => sig0000056a,
      C(37) => sig0000056a,
      C(36) => sig0000056a,
      C(35) => sig0000056a,
      C(34) => sig0000056a,
      C(33) => sig0000056a,
      C(32) => sig0000056a,
      C(31) => sig0000056a,
      C(30) => sig0000056a,
      C(29) => sig0000056a,
      C(28) => sig0000056a,
      C(27) => sig0000056a,
      C(26) => sig0000056b,
      C(25) => sig0000056c,
      C(24) => sig0000056d,
      C(23) => sig0000056e,
      C(22) => sig0000056f,
      C(21) => sig00000570,
      C(20) => sig00000571,
      C(19) => sig00000572,
      C(18) => sig00000573,
      C(17) => sig00000574,
      C(16) => sig00000575,
      C(15) => sig00000576,
      C(14) => sig00000577,
      C(13) => sig00000578,
      C(12) => sig00000579,
      C(11) => sig0000057a,
      C(10) => sig0000057b,
      C(9) => sig0000057c,
      C(8) => sig0000057d,
      C(7) => sig0000057e,
      C(6) => sig0000057f,
      C(5) => sig00000580,
      C(4) => sig00000581,
      C(3) => sig00000582,
      C(2) => sig00000583,
      C(1) => sig00000584,
      C(0) => sig00000585,
      CARRYINSEL(2) => sig000008b6,
      CARRYINSEL(1) => sig000008b6,
      CARRYINSEL(0) => sig000008b6,
      OPMODE(6) => sig000008b6,
      OPMODE(5) => sig000006d1,
      OPMODE(4) => sig000006d1,
      OPMODE(3) => sig000008b6,
      OPMODE(2) => sig000006d1,
      OPMODE(1) => sig000008b6,
      OPMODE(0) => sig000006d1,
      BCIN(17) => sig000008b6,
      BCIN(16) => sig000008b6,
      BCIN(15) => sig000008b6,
      BCIN(14) => sig000008b6,
      BCIN(13) => sig000008b6,
      BCIN(12) => sig000008b6,
      BCIN(11) => sig000008b6,
      BCIN(10) => sig000008b6,
      BCIN(9) => sig000008b6,
      BCIN(8) => sig000008b6,
      BCIN(7) => sig000008b6,
      BCIN(6) => sig000008b6,
      BCIN(5) => sig000008b6,
      BCIN(4) => sig000008b6,
      BCIN(3) => sig000008b6,
      BCIN(2) => sig000008b6,
      BCIN(1) => sig000008b6,
      BCIN(0) => sig000008b6,
      ALUMODE(3) => sig000008b6,
      ALUMODE(2) => sig000008b6,
      ALUMODE(1) => sig000008b6,
      ALUMODE(0) => sig000008b6,
      PCOUT(47) => NLW_blk00000655_PCOUT_47_UNCONNECTED,
      PCOUT(46) => NLW_blk00000655_PCOUT_46_UNCONNECTED,
      PCOUT(45) => NLW_blk00000655_PCOUT_45_UNCONNECTED,
      PCOUT(44) => NLW_blk00000655_PCOUT_44_UNCONNECTED,
      PCOUT(43) => NLW_blk00000655_PCOUT_43_UNCONNECTED,
      PCOUT(42) => NLW_blk00000655_PCOUT_42_UNCONNECTED,
      PCOUT(41) => NLW_blk00000655_PCOUT_41_UNCONNECTED,
      PCOUT(40) => NLW_blk00000655_PCOUT_40_UNCONNECTED,
      PCOUT(39) => NLW_blk00000655_PCOUT_39_UNCONNECTED,
      PCOUT(38) => NLW_blk00000655_PCOUT_38_UNCONNECTED,
      PCOUT(37) => NLW_blk00000655_PCOUT_37_UNCONNECTED,
      PCOUT(36) => NLW_blk00000655_PCOUT_36_UNCONNECTED,
      PCOUT(35) => NLW_blk00000655_PCOUT_35_UNCONNECTED,
      PCOUT(34) => NLW_blk00000655_PCOUT_34_UNCONNECTED,
      PCOUT(33) => NLW_blk00000655_PCOUT_33_UNCONNECTED,
      PCOUT(32) => NLW_blk00000655_PCOUT_32_UNCONNECTED,
      PCOUT(31) => NLW_blk00000655_PCOUT_31_UNCONNECTED,
      PCOUT(30) => NLW_blk00000655_PCOUT_30_UNCONNECTED,
      PCOUT(29) => NLW_blk00000655_PCOUT_29_UNCONNECTED,
      PCOUT(28) => NLW_blk00000655_PCOUT_28_UNCONNECTED,
      PCOUT(27) => NLW_blk00000655_PCOUT_27_UNCONNECTED,
      PCOUT(26) => NLW_blk00000655_PCOUT_26_UNCONNECTED,
      PCOUT(25) => NLW_blk00000655_PCOUT_25_UNCONNECTED,
      PCOUT(24) => NLW_blk00000655_PCOUT_24_UNCONNECTED,
      PCOUT(23) => NLW_blk00000655_PCOUT_23_UNCONNECTED,
      PCOUT(22) => NLW_blk00000655_PCOUT_22_UNCONNECTED,
      PCOUT(21) => NLW_blk00000655_PCOUT_21_UNCONNECTED,
      PCOUT(20) => NLW_blk00000655_PCOUT_20_UNCONNECTED,
      PCOUT(19) => NLW_blk00000655_PCOUT_19_UNCONNECTED,
      PCOUT(18) => NLW_blk00000655_PCOUT_18_UNCONNECTED,
      PCOUT(17) => NLW_blk00000655_PCOUT_17_UNCONNECTED,
      PCOUT(16) => NLW_blk00000655_PCOUT_16_UNCONNECTED,
      PCOUT(15) => NLW_blk00000655_PCOUT_15_UNCONNECTED,
      PCOUT(14) => NLW_blk00000655_PCOUT_14_UNCONNECTED,
      PCOUT(13) => NLW_blk00000655_PCOUT_13_UNCONNECTED,
      PCOUT(12) => NLW_blk00000655_PCOUT_12_UNCONNECTED,
      PCOUT(11) => NLW_blk00000655_PCOUT_11_UNCONNECTED,
      PCOUT(10) => NLW_blk00000655_PCOUT_10_UNCONNECTED,
      PCOUT(9) => NLW_blk00000655_PCOUT_9_UNCONNECTED,
      PCOUT(8) => NLW_blk00000655_PCOUT_8_UNCONNECTED,
      PCOUT(7) => NLW_blk00000655_PCOUT_7_UNCONNECTED,
      PCOUT(6) => NLW_blk00000655_PCOUT_6_UNCONNECTED,
      PCOUT(5) => NLW_blk00000655_PCOUT_5_UNCONNECTED,
      PCOUT(4) => NLW_blk00000655_PCOUT_4_UNCONNECTED,
      PCOUT(3) => NLW_blk00000655_PCOUT_3_UNCONNECTED,
      PCOUT(2) => NLW_blk00000655_PCOUT_2_UNCONNECTED,
      PCOUT(1) => NLW_blk00000655_PCOUT_1_UNCONNECTED,
      PCOUT(0) => NLW_blk00000655_PCOUT_0_UNCONNECTED,
      P(47) => NLW_blk00000655_P_47_UNCONNECTED,
      P(46) => NLW_blk00000655_P_46_UNCONNECTED,
      P(45) => NLW_blk00000655_P_45_UNCONNECTED,
      P(44) => NLW_blk00000655_P_44_UNCONNECTED,
      P(43) => NLW_blk00000655_P_43_UNCONNECTED,
      P(42) => sig00000505,
      P(41) => sig00000506,
      P(40) => sig00000507,
      P(39) => sig00000508,
      P(38) => sig00000509,
      P(37) => sig0000050a,
      P(36) => sig0000050b,
      P(35) => sig0000050c,
      P(34) => sig0000050d,
      P(33) => sig0000050e,
      P(32) => sig0000050f,
      P(31) => sig00000510,
      P(30) => sig00000511,
      P(29) => sig00000512,
      P(28) => sig00000513,
      P(27) => sig00000514,
      P(26) => sig00000515,
      P(25) => sig000001ff,
      P(24) => sig000001fe,
      P(23) => sig000001fd,
      P(22) => sig000001fc,
      P(21) => sig000001fb,
      P(20) => sig000001fa,
      P(19) => sig000001f9,
      P(18) => sig000001f8,
      P(17) => sig000001f7,
      P(16) => sig000001f6,
      P(15) => sig000001f5,
      P(14) => sig000001f4,
      P(13) => sig000001f3,
      P(12) => sig000001f2,
      P(11) => sig000001f1,
      P(10) => sig000001f0,
      P(9) => sig000001ef,
      P(8) => sig000001ee,
      P(7) => sig000001ed,
      P(6) => sig000001ec,
      P(5) => sig0000052a,
      P(4) => sig0000052b,
      P(3) => sig0000052c,
      P(2) => sig0000052d,
      P(1) => sig0000052e,
      P(0) => sig0000052f,
      BCOUT(17) => NLW_blk00000655_BCOUT_17_UNCONNECTED,
      BCOUT(16) => NLW_blk00000655_BCOUT_16_UNCONNECTED,
      BCOUT(15) => NLW_blk00000655_BCOUT_15_UNCONNECTED,
      BCOUT(14) => NLW_blk00000655_BCOUT_14_UNCONNECTED,
      BCOUT(13) => NLW_blk00000655_BCOUT_13_UNCONNECTED,
      BCOUT(12) => NLW_blk00000655_BCOUT_12_UNCONNECTED,
      BCOUT(11) => NLW_blk00000655_BCOUT_11_UNCONNECTED,
      BCOUT(10) => NLW_blk00000655_BCOUT_10_UNCONNECTED,
      BCOUT(9) => NLW_blk00000655_BCOUT_9_UNCONNECTED,
      BCOUT(8) => NLW_blk00000655_BCOUT_8_UNCONNECTED,
      BCOUT(7) => NLW_blk00000655_BCOUT_7_UNCONNECTED,
      BCOUT(6) => NLW_blk00000655_BCOUT_6_UNCONNECTED,
      BCOUT(5) => NLW_blk00000655_BCOUT_5_UNCONNECTED,
      BCOUT(4) => NLW_blk00000655_BCOUT_4_UNCONNECTED,
      BCOUT(3) => NLW_blk00000655_BCOUT_3_UNCONNECTED,
      BCOUT(2) => NLW_blk00000655_BCOUT_2_UNCONNECTED,
      BCOUT(1) => NLW_blk00000655_BCOUT_1_UNCONNECTED,
      BCOUT(0) => NLW_blk00000655_BCOUT_0_UNCONNECTED,
      ACIN(29) => sig000008b6,
      ACIN(28) => sig000008b6,
      ACIN(27) => sig000008b6,
      ACIN(26) => sig000008b6,
      ACIN(25) => sig000008b6,
      ACIN(24) => sig000008b6,
      ACIN(23) => sig000008b6,
      ACIN(22) => sig000008b6,
      ACIN(21) => sig000008b6,
      ACIN(20) => sig000008b6,
      ACIN(19) => sig000008b6,
      ACIN(18) => sig000008b6,
      ACIN(17) => sig000008b6,
      ACIN(16) => sig000008b6,
      ACIN(15) => sig000008b6,
      ACIN(14) => sig000008b6,
      ACIN(13) => sig000008b6,
      ACIN(12) => sig000008b6,
      ACIN(11) => sig000008b6,
      ACIN(10) => sig000008b6,
      ACIN(9) => sig000008b6,
      ACIN(8) => sig000008b6,
      ACIN(7) => sig000008b6,
      ACIN(6) => sig000008b6,
      ACIN(5) => sig000008b6,
      ACIN(4) => sig000008b6,
      ACIN(3) => sig000008b6,
      ACIN(2) => sig000008b6,
      ACIN(1) => sig000008b6,
      ACIN(0) => sig000008b6,
      ACOUT(29) => NLW_blk00000655_ACOUT_29_UNCONNECTED,
      ACOUT(28) => NLW_blk00000655_ACOUT_28_UNCONNECTED,
      ACOUT(27) => NLW_blk00000655_ACOUT_27_UNCONNECTED,
      ACOUT(26) => NLW_blk00000655_ACOUT_26_UNCONNECTED,
      ACOUT(25) => NLW_blk00000655_ACOUT_25_UNCONNECTED,
      ACOUT(24) => NLW_blk00000655_ACOUT_24_UNCONNECTED,
      ACOUT(23) => NLW_blk00000655_ACOUT_23_UNCONNECTED,
      ACOUT(22) => NLW_blk00000655_ACOUT_22_UNCONNECTED,
      ACOUT(21) => NLW_blk00000655_ACOUT_21_UNCONNECTED,
      ACOUT(20) => NLW_blk00000655_ACOUT_20_UNCONNECTED,
      ACOUT(19) => NLW_blk00000655_ACOUT_19_UNCONNECTED,
      ACOUT(18) => NLW_blk00000655_ACOUT_18_UNCONNECTED,
      ACOUT(17) => NLW_blk00000655_ACOUT_17_UNCONNECTED,
      ACOUT(16) => NLW_blk00000655_ACOUT_16_UNCONNECTED,
      ACOUT(15) => NLW_blk00000655_ACOUT_15_UNCONNECTED,
      ACOUT(14) => NLW_blk00000655_ACOUT_14_UNCONNECTED,
      ACOUT(13) => NLW_blk00000655_ACOUT_13_UNCONNECTED,
      ACOUT(12) => NLW_blk00000655_ACOUT_12_UNCONNECTED,
      ACOUT(11) => NLW_blk00000655_ACOUT_11_UNCONNECTED,
      ACOUT(10) => NLW_blk00000655_ACOUT_10_UNCONNECTED,
      ACOUT(9) => NLW_blk00000655_ACOUT_9_UNCONNECTED,
      ACOUT(8) => NLW_blk00000655_ACOUT_8_UNCONNECTED,
      ACOUT(7) => NLW_blk00000655_ACOUT_7_UNCONNECTED,
      ACOUT(6) => NLW_blk00000655_ACOUT_6_UNCONNECTED,
      ACOUT(5) => NLW_blk00000655_ACOUT_5_UNCONNECTED,
      ACOUT(4) => NLW_blk00000655_ACOUT_4_UNCONNECTED,
      ACOUT(3) => NLW_blk00000655_ACOUT_3_UNCONNECTED,
      ACOUT(2) => NLW_blk00000655_ACOUT_2_UNCONNECTED,
      ACOUT(1) => NLW_blk00000655_ACOUT_1_UNCONNECTED,
      ACOUT(0) => NLW_blk00000655_ACOUT_0_UNCONNECTED,
      CARRYOUT(3) => NLW_blk00000655_CARRYOUT_3_UNCONNECTED,
      CARRYOUT(2) => NLW_blk00000655_CARRYOUT_2_UNCONNECTED,
      CARRYOUT(1) => NLW_blk00000655_CARRYOUT_1_UNCONNECTED,
      CARRYOUT(0) => NLW_blk00000655_CARRYOUT_0_UNCONNECTED
    );
  blk00000656 : DSP48E
    generic map(
      ACASCREG => 2,
      ALUMODEREG => 0,
      AREG => 2,
      AUTORESET_PATTERN_DETECT => FALSE,
      AUTORESET_PATTERN_DETECT_OPTINV => "MATCH",
      A_INPUT => "DIRECT",
      BCASCREG => 1,
      BREG => 1,
      B_INPUT => "DIRECT",
      CARRYINREG => 0,
      CARRYINSELREG => 0,
      CREG => 0,
      MASK => X"000000000000",
      MREG => 1,
      MULTCARRYINREG => 0,
      OPMODEREG => 0,
      PATTERN => X"000000000000",
      PREG => 1,
      SEL_MASK => "MASK",
      SEL_PATTERN => "PATTERN",
      SEL_ROUNDING_MASK => "SEL_MASK",
      SIM_MODE => "SAFE",
      USE_MULT => "MULT_S",
      USE_PATTERN_DETECT => "NO_PATDET",
      USE_SIMD => "ONE48"
    )
    port map (
      CARRYIN => sig000008b6,
      CEA1 => ce,
      CEA2 => ce,
      CEB1 => sig000008b6,
      CEB2 => ce,
      CEC => sig000008b6,
      CECTRL => sig000008b6,
      CEP => ce,
      CEM => ce,
      CECARRYIN => sig000008b6,
      CEMULTCARRYIN => sig000008b6,
      CLK => clk,
      RSTA => sig000008b6,
      RSTB => sig000008b6,
      RSTC => sig000008b6,
      RSTCTRL => sig000008b6,
      RSTP => sig000008b6,
      RSTM => sig000008b6,
      RSTALLCARRYIN => sig000008b6,
      CEALUMODE => sig000008b6,
      RSTALUMODE => sig000008b6,
      PATTERNBDETECT => NLW_blk00000656_PATTERNBDETECT_UNCONNECTED,
      PATTERNDETECT => NLW_blk00000656_PATTERNDETECT_UNCONNECTED,
      OVERFLOW => NLW_blk00000656_OVERFLOW_UNCONNECTED,
      UNDERFLOW => NLW_blk00000656_UNDERFLOW_UNCONNECTED,
      CARRYCASCIN => sig000008b6,
      CARRYCASCOUT => NLW_blk00000656_CARRYCASCOUT_UNCONNECTED,
      MULTSIGNIN => sig000008b6,
      MULTSIGNOUT => NLW_blk00000656_MULTSIGNOUT_UNCONNECTED,
      A(29) => sig000008b6,
      A(28) => sig000008b6,
      A(27) => sig000008b6,
      A(26) => sig000008b6,
      A(25) => sig000008b6,
      A(24) => sig00000586,
      A(23) => sig00000586,
      A(22) => sig00000586,
      A(21) => sig00000586,
      A(20) => sig00000586,
      A(19) => sig00000586,
      A(18) => sig00000586,
      A(17) => sig00000586,
      A(16) => sig00000586,
      A(15) => sig00000586,
      A(14) => sig00000586,
      A(13) => sig00000586,
      A(12) => sig00000592,
      A(11) => sig00000593,
      A(10) => sig00000594,
      A(9) => sig00000595,
      A(8) => sig00000596,
      A(7) => sig00000597,
      A(6) => sig00000598,
      A(5) => sig00000599,
      A(4) => sig0000059a,
      A(3) => sig0000059b,
      A(2) => sig0000059c,
      A(1) => sig0000059d,
      A(0) => sig0000059e,
      PCIN(47) => sig000008b6,
      PCIN(46) => sig000008b6,
      PCIN(45) => sig000008b6,
      PCIN(44) => sig000008b6,
      PCIN(43) => sig000008b6,
      PCIN(42) => sig000008b6,
      PCIN(41) => sig000008b6,
      PCIN(40) => sig000008b6,
      PCIN(39) => sig000008b6,
      PCIN(38) => sig000008b6,
      PCIN(37) => sig000008b6,
      PCIN(36) => sig000008b6,
      PCIN(35) => sig000008b6,
      PCIN(34) => sig000008b6,
      PCIN(33) => sig000008b6,
      PCIN(32) => sig000008b6,
      PCIN(31) => sig000008b6,
      PCIN(30) => sig000008b6,
      PCIN(29) => sig000008b6,
      PCIN(28) => sig000008b6,
      PCIN(27) => sig000008b6,
      PCIN(26) => sig000008b6,
      PCIN(25) => sig000008b6,
      PCIN(24) => sig000008b6,
      PCIN(23) => sig000008b6,
      PCIN(22) => sig000008b6,
      PCIN(21) => sig000008b6,
      PCIN(20) => sig000008b6,
      PCIN(19) => sig000008b6,
      PCIN(18) => sig000008b6,
      PCIN(17) => sig000008b6,
      PCIN(16) => sig000008b6,
      PCIN(15) => sig000008b6,
      PCIN(14) => sig000008b6,
      PCIN(13) => sig000008b6,
      PCIN(12) => sig000008b6,
      PCIN(11) => sig000008b6,
      PCIN(10) => sig000008b6,
      PCIN(9) => sig000008b6,
      PCIN(8) => sig000008b6,
      PCIN(7) => sig000008b6,
      PCIN(6) => sig000008b6,
      PCIN(5) => sig000008b6,
      PCIN(4) => sig000008b6,
      PCIN(3) => sig000008b6,
      PCIN(2) => sig000008b6,
      PCIN(1) => sig000008b6,
      PCIN(0) => sig000008b6,
      B(17) => sig0000059f,
      B(16) => sig0000059f,
      B(15) => sig0000059f,
      B(14) => sig0000059f,
      B(13) => sig0000059f,
      B(12) => sig000005a4,
      B(11) => sig000005a5,
      B(10) => sig000005a6,
      B(9) => sig000005a7,
      B(8) => sig000005a8,
      B(7) => sig000005a9,
      B(6) => sig000005aa,
      B(5) => sig000005ab,
      B(4) => sig000005ac,
      B(3) => sig000005ad,
      B(2) => sig000005ae,
      B(1) => sig000005af,
      B(0) => sig000005b0,
      C(47) => sig000008b6,
      C(46) => sig000008b6,
      C(45) => sig000008b6,
      C(44) => sig000008b6,
      C(43) => sig000008b6,
      C(42) => sig000008b6,
      C(41) => sig000008b6,
      C(40) => sig000008b6,
      C(39) => sig000008b6,
      C(38) => sig000008b6,
      C(37) => sig000008b6,
      C(36) => sig000008b6,
      C(35) => sig000008b6,
      C(34) => sig000008b6,
      C(33) => sig000008b6,
      C(32) => sig000008b6,
      C(31) => sig000008b6,
      C(30) => sig000008b6,
      C(29) => sig000008b6,
      C(28) => sig000008b6,
      C(27) => sig000008b6,
      C(26) => sig000008b6,
      C(25) => sig000008b6,
      C(24) => sig000008b6,
      C(23) => sig000008b6,
      C(22) => sig000008b6,
      C(21) => sig000008b6,
      C(20) => sig000008b6,
      C(19) => sig000008b6,
      C(18) => sig000008b6,
      C(17) => sig000008b6,
      C(16) => sig000008b6,
      C(15) => sig000008b6,
      C(14) => sig000008b6,
      C(13) => sig000008b6,
      C(12) => sig000008b6,
      C(11) => sig000008b6,
      C(10) => sig000008b6,
      C(9) => sig000008b6,
      C(8) => sig000008b6,
      C(7) => sig000008b6,
      C(6) => sig000008b6,
      C(5) => sig000008b6,
      C(4) => sig000006d1,
      C(3) => sig000006d1,
      C(2) => sig000006d1,
      C(1) => sig000006d1,
      C(0) => sig000006d1,
      CARRYINSEL(2) => sig000008b6,
      CARRYINSEL(1) => sig000008b6,
      CARRYINSEL(0) => sig000008b6,
      OPMODE(6) => sig000008b6,
      OPMODE(5) => sig000006d1,
      OPMODE(4) => sig000006d1,
      OPMODE(3) => sig000008b6,
      OPMODE(2) => sig000006d1,
      OPMODE(1) => sig000008b6,
      OPMODE(0) => sig000006d1,
      BCIN(17) => sig000008b6,
      BCIN(16) => sig000008b6,
      BCIN(15) => sig000008b6,
      BCIN(14) => sig000008b6,
      BCIN(13) => sig000008b6,
      BCIN(12) => sig000008b6,
      BCIN(11) => sig000008b6,
      BCIN(10) => sig000008b6,
      BCIN(9) => sig000008b6,
      BCIN(8) => sig000008b6,
      BCIN(7) => sig000008b6,
      BCIN(6) => sig000008b6,
      BCIN(5) => sig000008b6,
      BCIN(4) => sig000008b6,
      BCIN(3) => sig000008b6,
      BCIN(2) => sig000008b6,
      BCIN(1) => sig000008b6,
      BCIN(0) => sig000008b6,
      ALUMODE(3) => sig000008b6,
      ALUMODE(2) => sig000008b6,
      ALUMODE(1) => sig000008b6,
      ALUMODE(0) => sig000008b6,
      PCOUT(47) => NLW_blk00000656_PCOUT_47_UNCONNECTED,
      PCOUT(46) => NLW_blk00000656_PCOUT_46_UNCONNECTED,
      PCOUT(45) => NLW_blk00000656_PCOUT_45_UNCONNECTED,
      PCOUT(44) => NLW_blk00000656_PCOUT_44_UNCONNECTED,
      PCOUT(43) => NLW_blk00000656_PCOUT_43_UNCONNECTED,
      PCOUT(42) => NLW_blk00000656_PCOUT_42_UNCONNECTED,
      PCOUT(41) => NLW_blk00000656_PCOUT_41_UNCONNECTED,
      PCOUT(40) => NLW_blk00000656_PCOUT_40_UNCONNECTED,
      PCOUT(39) => NLW_blk00000656_PCOUT_39_UNCONNECTED,
      PCOUT(38) => NLW_blk00000656_PCOUT_38_UNCONNECTED,
      PCOUT(37) => NLW_blk00000656_PCOUT_37_UNCONNECTED,
      PCOUT(36) => NLW_blk00000656_PCOUT_36_UNCONNECTED,
      PCOUT(35) => NLW_blk00000656_PCOUT_35_UNCONNECTED,
      PCOUT(34) => NLW_blk00000656_PCOUT_34_UNCONNECTED,
      PCOUT(33) => NLW_blk00000656_PCOUT_33_UNCONNECTED,
      PCOUT(32) => NLW_blk00000656_PCOUT_32_UNCONNECTED,
      PCOUT(31) => NLW_blk00000656_PCOUT_31_UNCONNECTED,
      PCOUT(30) => NLW_blk00000656_PCOUT_30_UNCONNECTED,
      PCOUT(29) => NLW_blk00000656_PCOUT_29_UNCONNECTED,
      PCOUT(28) => NLW_blk00000656_PCOUT_28_UNCONNECTED,
      PCOUT(27) => NLW_blk00000656_PCOUT_27_UNCONNECTED,
      PCOUT(26) => NLW_blk00000656_PCOUT_26_UNCONNECTED,
      PCOUT(25) => NLW_blk00000656_PCOUT_25_UNCONNECTED,
      PCOUT(24) => NLW_blk00000656_PCOUT_24_UNCONNECTED,
      PCOUT(23) => NLW_blk00000656_PCOUT_23_UNCONNECTED,
      PCOUT(22) => NLW_blk00000656_PCOUT_22_UNCONNECTED,
      PCOUT(21) => NLW_blk00000656_PCOUT_21_UNCONNECTED,
      PCOUT(20) => NLW_blk00000656_PCOUT_20_UNCONNECTED,
      PCOUT(19) => NLW_blk00000656_PCOUT_19_UNCONNECTED,
      PCOUT(18) => NLW_blk00000656_PCOUT_18_UNCONNECTED,
      PCOUT(17) => NLW_blk00000656_PCOUT_17_UNCONNECTED,
      PCOUT(16) => NLW_blk00000656_PCOUT_16_UNCONNECTED,
      PCOUT(15) => NLW_blk00000656_PCOUT_15_UNCONNECTED,
      PCOUT(14) => NLW_blk00000656_PCOUT_14_UNCONNECTED,
      PCOUT(13) => NLW_blk00000656_PCOUT_13_UNCONNECTED,
      PCOUT(12) => NLW_blk00000656_PCOUT_12_UNCONNECTED,
      PCOUT(11) => NLW_blk00000656_PCOUT_11_UNCONNECTED,
      PCOUT(10) => NLW_blk00000656_PCOUT_10_UNCONNECTED,
      PCOUT(9) => NLW_blk00000656_PCOUT_9_UNCONNECTED,
      PCOUT(8) => NLW_blk00000656_PCOUT_8_UNCONNECTED,
      PCOUT(7) => NLW_blk00000656_PCOUT_7_UNCONNECTED,
      PCOUT(6) => NLW_blk00000656_PCOUT_6_UNCONNECTED,
      PCOUT(5) => NLW_blk00000656_PCOUT_5_UNCONNECTED,
      PCOUT(4) => NLW_blk00000656_PCOUT_4_UNCONNECTED,
      PCOUT(3) => NLW_blk00000656_PCOUT_3_UNCONNECTED,
      PCOUT(2) => NLW_blk00000656_PCOUT_2_UNCONNECTED,
      PCOUT(1) => NLW_blk00000656_PCOUT_1_UNCONNECTED,
      PCOUT(0) => NLW_blk00000656_PCOUT_0_UNCONNECTED,
      P(47) => NLW_blk00000656_P_47_UNCONNECTED,
      P(46) => NLW_blk00000656_P_46_UNCONNECTED,
      P(45) => NLW_blk00000656_P_45_UNCONNECTED,
      P(44) => NLW_blk00000656_P_44_UNCONNECTED,
      P(43) => NLW_blk00000656_P_43_UNCONNECTED,
      P(42) => sig0000055b,
      P(41) => sig0000055c,
      P(40) => sig0000055d,
      P(39) => sig0000055e,
      P(38) => sig0000055f,
      P(37) => sig00000560,
      P(36) => sig00000561,
      P(35) => sig00000562,
      P(34) => sig00000563,
      P(33) => sig00000564,
      P(32) => sig00000565,
      P(31) => sig00000566,
      P(30) => sig00000567,
      P(29) => sig00000568,
      P(28) => sig00000569,
      P(27) => sig0000056a,
      P(26) => sig0000056b,
      P(25) => sig0000056c,
      P(24) => sig0000056d,
      P(23) => sig0000056e,
      P(22) => sig0000056f,
      P(21) => sig00000570,
      P(20) => sig00000571,
      P(19) => sig00000572,
      P(18) => sig00000573,
      P(17) => sig00000574,
      P(16) => sig00000575,
      P(15) => sig00000576,
      P(14) => sig00000577,
      P(13) => sig00000578,
      P(12) => sig00000579,
      P(11) => sig0000057a,
      P(10) => sig0000057b,
      P(9) => sig0000057c,
      P(8) => sig0000057d,
      P(7) => sig0000057e,
      P(6) => sig0000057f,
      P(5) => sig00000580,
      P(4) => sig00000581,
      P(3) => sig00000582,
      P(2) => sig00000583,
      P(1) => sig00000584,
      P(0) => sig00000585,
      BCOUT(17) => NLW_blk00000656_BCOUT_17_UNCONNECTED,
      BCOUT(16) => NLW_blk00000656_BCOUT_16_UNCONNECTED,
      BCOUT(15) => NLW_blk00000656_BCOUT_15_UNCONNECTED,
      BCOUT(14) => NLW_blk00000656_BCOUT_14_UNCONNECTED,
      BCOUT(13) => NLW_blk00000656_BCOUT_13_UNCONNECTED,
      BCOUT(12) => NLW_blk00000656_BCOUT_12_UNCONNECTED,
      BCOUT(11) => NLW_blk00000656_BCOUT_11_UNCONNECTED,
      BCOUT(10) => NLW_blk00000656_BCOUT_10_UNCONNECTED,
      BCOUT(9) => NLW_blk00000656_BCOUT_9_UNCONNECTED,
      BCOUT(8) => NLW_blk00000656_BCOUT_8_UNCONNECTED,
      BCOUT(7) => NLW_blk00000656_BCOUT_7_UNCONNECTED,
      BCOUT(6) => NLW_blk00000656_BCOUT_6_UNCONNECTED,
      BCOUT(5) => NLW_blk00000656_BCOUT_5_UNCONNECTED,
      BCOUT(4) => NLW_blk00000656_BCOUT_4_UNCONNECTED,
      BCOUT(3) => NLW_blk00000656_BCOUT_3_UNCONNECTED,
      BCOUT(2) => NLW_blk00000656_BCOUT_2_UNCONNECTED,
      BCOUT(1) => NLW_blk00000656_BCOUT_1_UNCONNECTED,
      BCOUT(0) => NLW_blk00000656_BCOUT_0_UNCONNECTED,
      ACIN(29) => sig000008b6,
      ACIN(28) => sig000008b6,
      ACIN(27) => sig000008b6,
      ACIN(26) => sig000008b6,
      ACIN(25) => sig000008b6,
      ACIN(24) => sig000008b6,
      ACIN(23) => sig000008b6,
      ACIN(22) => sig000008b6,
      ACIN(21) => sig000008b6,
      ACIN(20) => sig000008b6,
      ACIN(19) => sig000008b6,
      ACIN(18) => sig000008b6,
      ACIN(17) => sig000008b6,
      ACIN(16) => sig000008b6,
      ACIN(15) => sig000008b6,
      ACIN(14) => sig000008b6,
      ACIN(13) => sig000008b6,
      ACIN(12) => sig000008b6,
      ACIN(11) => sig000008b6,
      ACIN(10) => sig000008b6,
      ACIN(9) => sig000008b6,
      ACIN(8) => sig000008b6,
      ACIN(7) => sig000008b6,
      ACIN(6) => sig000008b6,
      ACIN(5) => sig000008b6,
      ACIN(4) => sig000008b6,
      ACIN(3) => sig000008b6,
      ACIN(2) => sig000008b6,
      ACIN(1) => sig000008b6,
      ACIN(0) => sig000008b6,
      ACOUT(29) => NLW_blk00000656_ACOUT_29_UNCONNECTED,
      ACOUT(28) => NLW_blk00000656_ACOUT_28_UNCONNECTED,
      ACOUT(27) => NLW_blk00000656_ACOUT_27_UNCONNECTED,
      ACOUT(26) => NLW_blk00000656_ACOUT_26_UNCONNECTED,
      ACOUT(25) => NLW_blk00000656_ACOUT_25_UNCONNECTED,
      ACOUT(24) => NLW_blk00000656_ACOUT_24_UNCONNECTED,
      ACOUT(23) => NLW_blk00000656_ACOUT_23_UNCONNECTED,
      ACOUT(22) => NLW_blk00000656_ACOUT_22_UNCONNECTED,
      ACOUT(21) => NLW_blk00000656_ACOUT_21_UNCONNECTED,
      ACOUT(20) => NLW_blk00000656_ACOUT_20_UNCONNECTED,
      ACOUT(19) => NLW_blk00000656_ACOUT_19_UNCONNECTED,
      ACOUT(18) => NLW_blk00000656_ACOUT_18_UNCONNECTED,
      ACOUT(17) => NLW_blk00000656_ACOUT_17_UNCONNECTED,
      ACOUT(16) => NLW_blk00000656_ACOUT_16_UNCONNECTED,
      ACOUT(15) => NLW_blk00000656_ACOUT_15_UNCONNECTED,
      ACOUT(14) => NLW_blk00000656_ACOUT_14_UNCONNECTED,
      ACOUT(13) => NLW_blk00000656_ACOUT_13_UNCONNECTED,
      ACOUT(12) => NLW_blk00000656_ACOUT_12_UNCONNECTED,
      ACOUT(11) => NLW_blk00000656_ACOUT_11_UNCONNECTED,
      ACOUT(10) => NLW_blk00000656_ACOUT_10_UNCONNECTED,
      ACOUT(9) => NLW_blk00000656_ACOUT_9_UNCONNECTED,
      ACOUT(8) => NLW_blk00000656_ACOUT_8_UNCONNECTED,
      ACOUT(7) => NLW_blk00000656_ACOUT_7_UNCONNECTED,
      ACOUT(6) => NLW_blk00000656_ACOUT_6_UNCONNECTED,
      ACOUT(5) => NLW_blk00000656_ACOUT_5_UNCONNECTED,
      ACOUT(4) => NLW_blk00000656_ACOUT_4_UNCONNECTED,
      ACOUT(3) => NLW_blk00000656_ACOUT_3_UNCONNECTED,
      ACOUT(2) => NLW_blk00000656_ACOUT_2_UNCONNECTED,
      ACOUT(1) => NLW_blk00000656_ACOUT_1_UNCONNECTED,
      ACOUT(0) => NLW_blk00000656_ACOUT_0_UNCONNECTED,
      CARRYOUT(3) => NLW_blk00000656_CARRYOUT_3_UNCONNECTED,
      CARRYOUT(2) => NLW_blk00000656_CARRYOUT_2_UNCONNECTED,
      CARRYOUT(1) => NLW_blk00000656_CARRYOUT_1_UNCONNECTED,
      CARRYOUT(0) => NLW_blk00000656_CARRYOUT_0_UNCONNECTED
    );
  blk00000657 : DSP48E
    generic map(
      ACASCREG => 2,
      ALUMODEREG => 0,
      AREG => 2,
      AUTORESET_PATTERN_DETECT => FALSE,
      AUTORESET_PATTERN_DETECT_OPTINV => "MATCH",
      A_INPUT => "DIRECT",
      BCASCREG => 2,
      BREG => 2,
      B_INPUT => "DIRECT",
      CARRYINREG => 0,
      CARRYINSELREG => 0,
      CREG => 1,
      MASK => X"000000000000",
      MREG => 1,
      MULTCARRYINREG => 0,
      OPMODEREG => 0,
      PATTERN => X"000000000000",
      PREG => 1,
      SEL_MASK => "MASK",
      SEL_PATTERN => "PATTERN",
      SEL_ROUNDING_MASK => "SEL_MASK",
      SIM_MODE => "SAFE",
      USE_MULT => "MULT_S",
      USE_PATTERN_DETECT => "NO_PATDET",
      USE_SIMD => "ONE48"
    )
    port map (
      CARRYIN => sig000008b6,
      CEA1 => ce,
      CEA2 => ce,
      CEB1 => ce,
      CEB2 => ce,
      CEC => ce,
      CECTRL => sig000008b6,
      CEP => ce,
      CEM => ce,
      CECARRYIN => sig000008b6,
      CEMULTCARRYIN => sig000008b6,
      CLK => clk,
      RSTA => sig000008b6,
      RSTB => sig000008b6,
      RSTC => sig000008b6,
      RSTCTRL => sig000008b6,
      RSTP => sig000008b6,
      RSTM => sig000008b6,
      RSTALLCARRYIN => sig000008b6,
      CEALUMODE => sig000008b6,
      RSTALUMODE => sig000008b6,
      PATTERNBDETECT => NLW_blk00000657_PATTERNBDETECT_UNCONNECTED,
      PATTERNDETECT => NLW_blk00000657_PATTERNDETECT_UNCONNECTED,
      OVERFLOW => NLW_blk00000657_OVERFLOW_UNCONNECTED,
      UNDERFLOW => NLW_blk00000657_UNDERFLOW_UNCONNECTED,
      CARRYCASCIN => sig000008b6,
      CARRYCASCOUT => NLW_blk00000657_CARRYCASCOUT_UNCONNECTED,
      MULTSIGNIN => sig000008b6,
      MULTSIGNOUT => NLW_blk00000657_MULTSIGNOUT_UNCONNECTED,
      A(29) => sig000008b6,
      A(28) => sig000008b6,
      A(27) => sig000008b6,
      A(26) => sig000008b6,
      A(25) => sig000008b6,
      A(24) => sig000005dc,
      A(23) => sig000005dc,
      A(22) => sig000005dc,
      A(21) => sig000005dc,
      A(20) => sig000005dc,
      A(19) => sig000005dc,
      A(18) => sig000005dc,
      A(17) => sig000005dc,
      A(16) => sig000005dc,
      A(15) => sig000005dc,
      A(14) => sig000005dc,
      A(13) => sig000005dc,
      A(12) => sig000005dc,
      A(11) => sig000005e9,
      A(10) => sig000005ea,
      A(9) => sig000005eb,
      A(8) => sig000005ec,
      A(7) => sig000005ed,
      A(6) => sig000005ee,
      A(5) => sig000005ef,
      A(4) => sig000005f0,
      A(3) => sig000005f1,
      A(2) => sig000005f2,
      A(1) => sig000005f3,
      A(0) => sig000005f4,
      PCIN(47) => sig000008b6,
      PCIN(46) => sig000008b6,
      PCIN(45) => sig000008b6,
      PCIN(44) => sig000008b6,
      PCIN(43) => sig000008b6,
      PCIN(42) => sig000008b6,
      PCIN(41) => sig000008b6,
      PCIN(40) => sig000008b6,
      PCIN(39) => sig000008b6,
      PCIN(38) => sig000008b6,
      PCIN(37) => sig000008b6,
      PCIN(36) => sig000008b6,
      PCIN(35) => sig000008b6,
      PCIN(34) => sig000008b6,
      PCIN(33) => sig000008b6,
      PCIN(32) => sig000008b6,
      PCIN(31) => sig000008b6,
      PCIN(30) => sig000008b6,
      PCIN(29) => sig000008b6,
      PCIN(28) => sig000008b6,
      PCIN(27) => sig000008b6,
      PCIN(26) => sig000008b6,
      PCIN(25) => sig000008b6,
      PCIN(24) => sig000008b6,
      PCIN(23) => sig000008b6,
      PCIN(22) => sig000008b6,
      PCIN(21) => sig000008b6,
      PCIN(20) => sig000008b6,
      PCIN(19) => sig000008b6,
      PCIN(18) => sig000008b6,
      PCIN(17) => sig000008b6,
      PCIN(16) => sig000008b6,
      PCIN(15) => sig000008b6,
      PCIN(14) => sig000008b6,
      PCIN(13) => sig000008b6,
      PCIN(12) => sig000008b6,
      PCIN(11) => sig000008b6,
      PCIN(10) => sig000008b6,
      PCIN(9) => sig000008b6,
      PCIN(8) => sig000008b6,
      PCIN(7) => sig000008b6,
      PCIN(6) => sig000008b6,
      PCIN(5) => sig000008b6,
      PCIN(4) => sig000008b6,
      PCIN(3) => sig000008b6,
      PCIN(2) => sig000008b6,
      PCIN(1) => sig000008b6,
      PCIN(0) => sig000008b6,
      B(17) => sig000005f5,
      B(16) => sig000005f5,
      B(15) => sig000005f5,
      B(14) => sig000005f5,
      B(13) => sig000005f9,
      B(12) => sig000005fa,
      B(11) => sig000005fb,
      B(10) => sig000005fc,
      B(9) => sig000005fd,
      B(8) => sig000005fe,
      B(7) => sig000005ff,
      B(6) => sig00000600,
      B(5) => sig00000601,
      B(4) => sig00000602,
      B(3) => sig00000603,
      B(2) => sig00000604,
      B(1) => sig00000605,
      B(0) => sig0000055a,
      C(47) => sig0000056a,
      C(46) => sig0000056a,
      C(45) => sig0000056a,
      C(44) => sig0000056a,
      C(43) => sig0000056a,
      C(42) => sig0000056a,
      C(41) => sig0000056a,
      C(40) => sig0000056a,
      C(39) => sig0000056a,
      C(38) => sig0000056a,
      C(37) => sig0000056a,
      C(36) => sig0000056a,
      C(35) => sig0000056a,
      C(34) => sig0000056a,
      C(33) => sig0000056a,
      C(32) => sig0000056a,
      C(31) => sig0000056a,
      C(30) => sig0000056a,
      C(29) => sig0000056a,
      C(28) => sig0000056a,
      C(27) => sig0000056a,
      C(26) => sig0000056b,
      C(25) => sig0000056c,
      C(24) => sig0000056d,
      C(23) => sig0000056e,
      C(22) => sig0000056f,
      C(21) => sig00000570,
      C(20) => sig00000571,
      C(19) => sig00000572,
      C(18) => sig00000573,
      C(17) => sig00000574,
      C(16) => sig00000575,
      C(15) => sig00000576,
      C(14) => sig00000577,
      C(13) => sig00000578,
      C(12) => sig00000579,
      C(11) => sig0000057a,
      C(10) => sig0000057b,
      C(9) => sig0000057c,
      C(8) => sig0000057d,
      C(7) => sig0000057e,
      C(6) => sig0000057f,
      C(5) => sig00000580,
      C(4) => sig00000581,
      C(3) => sig00000582,
      C(2) => sig00000583,
      C(1) => sig00000584,
      C(0) => sig00000585,
      CARRYINSEL(2) => sig000008b6,
      CARRYINSEL(1) => sig000008b6,
      CARRYINSEL(0) => sig000008b6,
      OPMODE(6) => sig000008b6,
      OPMODE(5) => sig000006d1,
      OPMODE(4) => sig000006d1,
      OPMODE(3) => sig000008b6,
      OPMODE(2) => sig000006d1,
      OPMODE(1) => sig000008b6,
      OPMODE(0) => sig000006d1,
      BCIN(17) => sig000008b6,
      BCIN(16) => sig000008b6,
      BCIN(15) => sig000008b6,
      BCIN(14) => sig000008b6,
      BCIN(13) => sig000008b6,
      BCIN(12) => sig000008b6,
      BCIN(11) => sig000008b6,
      BCIN(10) => sig000008b6,
      BCIN(9) => sig000008b6,
      BCIN(8) => sig000008b6,
      BCIN(7) => sig000008b6,
      BCIN(6) => sig000008b6,
      BCIN(5) => sig000008b6,
      BCIN(4) => sig000008b6,
      BCIN(3) => sig000008b6,
      BCIN(2) => sig000008b6,
      BCIN(1) => sig000008b6,
      BCIN(0) => sig000008b6,
      ALUMODE(3) => sig000008b6,
      ALUMODE(2) => sig000008b6,
      ALUMODE(1) => sig000006d1,
      ALUMODE(0) => sig000006d1,
      PCOUT(47) => NLW_blk00000657_PCOUT_47_UNCONNECTED,
      PCOUT(46) => NLW_blk00000657_PCOUT_46_UNCONNECTED,
      PCOUT(45) => NLW_blk00000657_PCOUT_45_UNCONNECTED,
      PCOUT(44) => NLW_blk00000657_PCOUT_44_UNCONNECTED,
      PCOUT(43) => NLW_blk00000657_PCOUT_43_UNCONNECTED,
      PCOUT(42) => NLW_blk00000657_PCOUT_42_UNCONNECTED,
      PCOUT(41) => NLW_blk00000657_PCOUT_41_UNCONNECTED,
      PCOUT(40) => NLW_blk00000657_PCOUT_40_UNCONNECTED,
      PCOUT(39) => NLW_blk00000657_PCOUT_39_UNCONNECTED,
      PCOUT(38) => NLW_blk00000657_PCOUT_38_UNCONNECTED,
      PCOUT(37) => NLW_blk00000657_PCOUT_37_UNCONNECTED,
      PCOUT(36) => NLW_blk00000657_PCOUT_36_UNCONNECTED,
      PCOUT(35) => NLW_blk00000657_PCOUT_35_UNCONNECTED,
      PCOUT(34) => NLW_blk00000657_PCOUT_34_UNCONNECTED,
      PCOUT(33) => NLW_blk00000657_PCOUT_33_UNCONNECTED,
      PCOUT(32) => NLW_blk00000657_PCOUT_32_UNCONNECTED,
      PCOUT(31) => NLW_blk00000657_PCOUT_31_UNCONNECTED,
      PCOUT(30) => NLW_blk00000657_PCOUT_30_UNCONNECTED,
      PCOUT(29) => NLW_blk00000657_PCOUT_29_UNCONNECTED,
      PCOUT(28) => NLW_blk00000657_PCOUT_28_UNCONNECTED,
      PCOUT(27) => NLW_blk00000657_PCOUT_27_UNCONNECTED,
      PCOUT(26) => NLW_blk00000657_PCOUT_26_UNCONNECTED,
      PCOUT(25) => NLW_blk00000657_PCOUT_25_UNCONNECTED,
      PCOUT(24) => NLW_blk00000657_PCOUT_24_UNCONNECTED,
      PCOUT(23) => NLW_blk00000657_PCOUT_23_UNCONNECTED,
      PCOUT(22) => NLW_blk00000657_PCOUT_22_UNCONNECTED,
      PCOUT(21) => NLW_blk00000657_PCOUT_21_UNCONNECTED,
      PCOUT(20) => NLW_blk00000657_PCOUT_20_UNCONNECTED,
      PCOUT(19) => NLW_blk00000657_PCOUT_19_UNCONNECTED,
      PCOUT(18) => NLW_blk00000657_PCOUT_18_UNCONNECTED,
      PCOUT(17) => NLW_blk00000657_PCOUT_17_UNCONNECTED,
      PCOUT(16) => NLW_blk00000657_PCOUT_16_UNCONNECTED,
      PCOUT(15) => NLW_blk00000657_PCOUT_15_UNCONNECTED,
      PCOUT(14) => NLW_blk00000657_PCOUT_14_UNCONNECTED,
      PCOUT(13) => NLW_blk00000657_PCOUT_13_UNCONNECTED,
      PCOUT(12) => NLW_blk00000657_PCOUT_12_UNCONNECTED,
      PCOUT(11) => NLW_blk00000657_PCOUT_11_UNCONNECTED,
      PCOUT(10) => NLW_blk00000657_PCOUT_10_UNCONNECTED,
      PCOUT(9) => NLW_blk00000657_PCOUT_9_UNCONNECTED,
      PCOUT(8) => NLW_blk00000657_PCOUT_8_UNCONNECTED,
      PCOUT(7) => NLW_blk00000657_PCOUT_7_UNCONNECTED,
      PCOUT(6) => NLW_blk00000657_PCOUT_6_UNCONNECTED,
      PCOUT(5) => NLW_blk00000657_PCOUT_5_UNCONNECTED,
      PCOUT(4) => NLW_blk00000657_PCOUT_4_UNCONNECTED,
      PCOUT(3) => NLW_blk00000657_PCOUT_3_UNCONNECTED,
      PCOUT(2) => NLW_blk00000657_PCOUT_2_UNCONNECTED,
      PCOUT(1) => NLW_blk00000657_PCOUT_1_UNCONNECTED,
      PCOUT(0) => NLW_blk00000657_PCOUT_0_UNCONNECTED,
      P(47) => NLW_blk00000657_P_47_UNCONNECTED,
      P(46) => NLW_blk00000657_P_46_UNCONNECTED,
      P(45) => NLW_blk00000657_P_45_UNCONNECTED,
      P(44) => NLW_blk00000657_P_44_UNCONNECTED,
      P(43) => NLW_blk00000657_P_43_UNCONNECTED,
      P(42) => sig000005b1,
      P(41) => sig000005b2,
      P(40) => sig000005b3,
      P(39) => sig000005b4,
      P(38) => sig000005b5,
      P(37) => sig000005b6,
      P(36) => sig000005b7,
      P(35) => sig000005b8,
      P(34) => sig000005b9,
      P(33) => sig000005ba,
      P(32) => sig000005bb,
      P(31) => sig000005bc,
      P(30) => sig000005bd,
      P(29) => sig000005be,
      P(28) => sig000005bf,
      P(27) => sig000005c0,
      P(26) => sig000005c1,
      P(25) => sig00000213,
      P(24) => sig00000212,
      P(23) => sig00000211,
      P(22) => sig00000210,
      P(21) => sig0000020f,
      P(20) => sig0000020e,
      P(19) => sig0000020d,
      P(18) => sig0000020c,
      P(17) => sig0000020b,
      P(16) => sig0000020a,
      P(15) => sig00000209,
      P(14) => sig00000208,
      P(13) => sig00000207,
      P(12) => sig00000206,
      P(11) => sig00000205,
      P(10) => sig00000204,
      P(9) => sig00000203,
      P(8) => sig00000202,
      P(7) => sig00000201,
      P(6) => sig00000200,
      P(5) => sig000005d6,
      P(4) => sig000005d7,
      P(3) => sig000005d8,
      P(2) => sig000005d9,
      P(1) => sig000005da,
      P(0) => sig000005db,
      BCOUT(17) => NLW_blk00000657_BCOUT_17_UNCONNECTED,
      BCOUT(16) => NLW_blk00000657_BCOUT_16_UNCONNECTED,
      BCOUT(15) => NLW_blk00000657_BCOUT_15_UNCONNECTED,
      BCOUT(14) => NLW_blk00000657_BCOUT_14_UNCONNECTED,
      BCOUT(13) => NLW_blk00000657_BCOUT_13_UNCONNECTED,
      BCOUT(12) => NLW_blk00000657_BCOUT_12_UNCONNECTED,
      BCOUT(11) => NLW_blk00000657_BCOUT_11_UNCONNECTED,
      BCOUT(10) => NLW_blk00000657_BCOUT_10_UNCONNECTED,
      BCOUT(9) => NLW_blk00000657_BCOUT_9_UNCONNECTED,
      BCOUT(8) => NLW_blk00000657_BCOUT_8_UNCONNECTED,
      BCOUT(7) => NLW_blk00000657_BCOUT_7_UNCONNECTED,
      BCOUT(6) => NLW_blk00000657_BCOUT_6_UNCONNECTED,
      BCOUT(5) => NLW_blk00000657_BCOUT_5_UNCONNECTED,
      BCOUT(4) => NLW_blk00000657_BCOUT_4_UNCONNECTED,
      BCOUT(3) => NLW_blk00000657_BCOUT_3_UNCONNECTED,
      BCOUT(2) => NLW_blk00000657_BCOUT_2_UNCONNECTED,
      BCOUT(1) => NLW_blk00000657_BCOUT_1_UNCONNECTED,
      BCOUT(0) => NLW_blk00000657_BCOUT_0_UNCONNECTED,
      ACIN(29) => sig000008b6,
      ACIN(28) => sig000008b6,
      ACIN(27) => sig000008b6,
      ACIN(26) => sig000008b6,
      ACIN(25) => sig000008b6,
      ACIN(24) => sig000008b6,
      ACIN(23) => sig000008b6,
      ACIN(22) => sig000008b6,
      ACIN(21) => sig000008b6,
      ACIN(20) => sig000008b6,
      ACIN(19) => sig000008b6,
      ACIN(18) => sig000008b6,
      ACIN(17) => sig000008b6,
      ACIN(16) => sig000008b6,
      ACIN(15) => sig000008b6,
      ACIN(14) => sig000008b6,
      ACIN(13) => sig000008b6,
      ACIN(12) => sig000008b6,
      ACIN(11) => sig000008b6,
      ACIN(10) => sig000008b6,
      ACIN(9) => sig000008b6,
      ACIN(8) => sig000008b6,
      ACIN(7) => sig000008b6,
      ACIN(6) => sig000008b6,
      ACIN(5) => sig000008b6,
      ACIN(4) => sig000008b6,
      ACIN(3) => sig000008b6,
      ACIN(2) => sig000008b6,
      ACIN(1) => sig000008b6,
      ACIN(0) => sig000008b6,
      ACOUT(29) => NLW_blk00000657_ACOUT_29_UNCONNECTED,
      ACOUT(28) => NLW_blk00000657_ACOUT_28_UNCONNECTED,
      ACOUT(27) => NLW_blk00000657_ACOUT_27_UNCONNECTED,
      ACOUT(26) => NLW_blk00000657_ACOUT_26_UNCONNECTED,
      ACOUT(25) => NLW_blk00000657_ACOUT_25_UNCONNECTED,
      ACOUT(24) => NLW_blk00000657_ACOUT_24_UNCONNECTED,
      ACOUT(23) => NLW_blk00000657_ACOUT_23_UNCONNECTED,
      ACOUT(22) => NLW_blk00000657_ACOUT_22_UNCONNECTED,
      ACOUT(21) => NLW_blk00000657_ACOUT_21_UNCONNECTED,
      ACOUT(20) => NLW_blk00000657_ACOUT_20_UNCONNECTED,
      ACOUT(19) => NLW_blk00000657_ACOUT_19_UNCONNECTED,
      ACOUT(18) => NLW_blk00000657_ACOUT_18_UNCONNECTED,
      ACOUT(17) => NLW_blk00000657_ACOUT_17_UNCONNECTED,
      ACOUT(16) => NLW_blk00000657_ACOUT_16_UNCONNECTED,
      ACOUT(15) => NLW_blk00000657_ACOUT_15_UNCONNECTED,
      ACOUT(14) => NLW_blk00000657_ACOUT_14_UNCONNECTED,
      ACOUT(13) => NLW_blk00000657_ACOUT_13_UNCONNECTED,
      ACOUT(12) => NLW_blk00000657_ACOUT_12_UNCONNECTED,
      ACOUT(11) => NLW_blk00000657_ACOUT_11_UNCONNECTED,
      ACOUT(10) => NLW_blk00000657_ACOUT_10_UNCONNECTED,
      ACOUT(9) => NLW_blk00000657_ACOUT_9_UNCONNECTED,
      ACOUT(8) => NLW_blk00000657_ACOUT_8_UNCONNECTED,
      ACOUT(7) => NLW_blk00000657_ACOUT_7_UNCONNECTED,
      ACOUT(6) => NLW_blk00000657_ACOUT_6_UNCONNECTED,
      ACOUT(5) => NLW_blk00000657_ACOUT_5_UNCONNECTED,
      ACOUT(4) => NLW_blk00000657_ACOUT_4_UNCONNECTED,
      ACOUT(3) => NLW_blk00000657_ACOUT_3_UNCONNECTED,
      ACOUT(2) => NLW_blk00000657_ACOUT_2_UNCONNECTED,
      ACOUT(1) => NLW_blk00000657_ACOUT_1_UNCONNECTED,
      ACOUT(0) => NLW_blk00000657_ACOUT_0_UNCONNECTED,
      CARRYOUT(3) => NLW_blk00000657_CARRYOUT_3_UNCONNECTED,
      CARRYOUT(2) => NLW_blk00000657_CARRYOUT_2_UNCONNECTED,
      CARRYOUT(1) => NLW_blk00000657_CARRYOUT_1_UNCONNECTED,
      CARRYOUT(0) => NLW_blk00000657_CARRYOUT_0_UNCONNECTED
    );
  blk00000658 : XORCY
    port map (
      CI => sig000004b1,
      LI => sig000004b0,
      O => sig00000622
    );
  blk00000659 : LUT2
    generic map(
      INIT => X"9"
    )
    port map (
      I0 => sig000006d0,
      I1 => sig00000586,
      O => sig000004b0
    );
  blk0000065a : XORCY
    port map (
      CI => sig000004b3,
      LI => sig000004b2,
      O => sig00000621
    );
  blk0000065b : MUXCY
    port map (
      CI => sig000004b3,
      DI => sig000006d0,
      S => sig000004b2,
      O => sig000004b1
    );
  blk0000065c : LUT2
    generic map(
      INIT => X"9"
    )
    port map (
      I0 => sig000006d0,
      I1 => sig00000586,
      O => sig000004b2
    );
  blk0000065d : XORCY
    port map (
      CI => sig000004b5,
      LI => sig000004b4,
      O => sig00000620
    );
  blk0000065e : MUXCY
    port map (
      CI => sig000004b5,
      DI => sig000006cf,
      S => sig000004b4,
      O => sig000004b3
    );
  blk0000065f : LUT2
    generic map(
      INIT => X"9"
    )
    port map (
      I0 => sig000006cf,
      I1 => sig00000592,
      O => sig000004b4
    );
  blk00000660 : XORCY
    port map (
      CI => sig000004b7,
      LI => sig000004b6,
      O => sig0000061f
    );
  blk00000661 : MUXCY
    port map (
      CI => sig000004b7,
      DI => sig000006ce,
      S => sig000004b6,
      O => sig000004b5
    );
  blk00000662 : LUT2
    generic map(
      INIT => X"9"
    )
    port map (
      I0 => sig000006ce,
      I1 => sig00000593,
      O => sig000004b6
    );
  blk00000663 : XORCY
    port map (
      CI => sig000004b9,
      LI => sig000004b8,
      O => sig0000061e
    );
  blk00000664 : MUXCY
    port map (
      CI => sig000004b9,
      DI => sig000006cd,
      S => sig000004b8,
      O => sig000004b7
    );
  blk00000665 : LUT2
    generic map(
      INIT => X"9"
    )
    port map (
      I0 => sig000006cd,
      I1 => sig00000594,
      O => sig000004b8
    );
  blk00000666 : XORCY
    port map (
      CI => sig000004bb,
      LI => sig000004ba,
      O => sig0000061d
    );
  blk00000667 : MUXCY
    port map (
      CI => sig000004bb,
      DI => sig000006cc,
      S => sig000004ba,
      O => sig000004b9
    );
  blk00000668 : LUT2
    generic map(
      INIT => X"9"
    )
    port map (
      I0 => sig000006cc,
      I1 => sig00000595,
      O => sig000004ba
    );
  blk00000669 : XORCY
    port map (
      CI => sig000004bd,
      LI => sig000004bc,
      O => sig0000061c
    );
  blk0000066a : MUXCY
    port map (
      CI => sig000004bd,
      DI => sig000006cb,
      S => sig000004bc,
      O => sig000004bb
    );
  blk0000066b : LUT2
    generic map(
      INIT => X"9"
    )
    port map (
      I0 => sig000006cb,
      I1 => sig00000596,
      O => sig000004bc
    );
  blk0000066c : XORCY
    port map (
      CI => sig000004bf,
      LI => sig000004be,
      O => sig0000061b
    );
  blk0000066d : MUXCY
    port map (
      CI => sig000004bf,
      DI => sig000006ca,
      S => sig000004be,
      O => sig000004bd
    );
  blk0000066e : LUT2
    generic map(
      INIT => X"9"
    )
    port map (
      I0 => sig000006ca,
      I1 => sig00000597,
      O => sig000004be
    );
  blk0000066f : XORCY
    port map (
      CI => sig000004c1,
      LI => sig000004c0,
      O => sig0000061a
    );
  blk00000670 : MUXCY
    port map (
      CI => sig000004c1,
      DI => sig000006c9,
      S => sig000004c0,
      O => sig000004bf
    );
  blk00000671 : LUT2
    generic map(
      INIT => X"9"
    )
    port map (
      I0 => sig000006c9,
      I1 => sig00000598,
      O => sig000004c0
    );
  blk00000672 : XORCY
    port map (
      CI => sig000004c3,
      LI => sig000004c2,
      O => sig00000619
    );
  blk00000673 : MUXCY
    port map (
      CI => sig000004c3,
      DI => sig000006c8,
      S => sig000004c2,
      O => sig000004c1
    );
  blk00000674 : LUT2
    generic map(
      INIT => X"9"
    )
    port map (
      I0 => sig000006c8,
      I1 => sig00000599,
      O => sig000004c2
    );
  blk00000675 : XORCY
    port map (
      CI => sig000004c5,
      LI => sig000004c4,
      O => sig00000618
    );
  blk00000676 : MUXCY
    port map (
      CI => sig000004c5,
      DI => sig000006c7,
      S => sig000004c4,
      O => sig000004c3
    );
  blk00000677 : LUT2
    generic map(
      INIT => X"9"
    )
    port map (
      I0 => sig000006c7,
      I1 => sig0000059a,
      O => sig000004c4
    );
  blk00000678 : XORCY
    port map (
      CI => sig000004c7,
      LI => sig000004c6,
      O => sig00000617
    );
  blk00000679 : MUXCY
    port map (
      CI => sig000004c7,
      DI => sig000006c6,
      S => sig000004c6,
      O => sig000004c5
    );
  blk0000067a : LUT2
    generic map(
      INIT => X"9"
    )
    port map (
      I0 => sig000006c6,
      I1 => sig0000059b,
      O => sig000004c6
    );
  blk0000067b : XORCY
    port map (
      CI => sig000004c9,
      LI => sig000004c8,
      O => sig00000616
    );
  blk0000067c : MUXCY
    port map (
      CI => sig000004c9,
      DI => sig000006c5,
      S => sig000004c8,
      O => sig000004c7
    );
  blk0000067d : LUT2
    generic map(
      INIT => X"9"
    )
    port map (
      I0 => sig000006c5,
      I1 => sig0000059c,
      O => sig000004c8
    );
  blk0000067e : XORCY
    port map (
      CI => sig000004cb,
      LI => sig000004ca,
      O => sig00000615
    );
  blk0000067f : MUXCY
    port map (
      CI => sig000004cb,
      DI => sig000006c4,
      S => sig000004ca,
      O => sig000004c9
    );
  blk00000680 : LUT2
    generic map(
      INIT => X"9"
    )
    port map (
      I0 => sig000006c4,
      I1 => sig0000059d,
      O => sig000004ca
    );
  blk00000681 : MUXCY
    port map (
      CI => sig000006d1,
      DI => sig000006c3,
      S => sig000004cc,
      O => sig000004cb
    );
  blk00000682 : LUT2
    generic map(
      INIT => X"9"
    )
    port map (
      I0 => sig000006c3,
      I1 => sig0000059e,
      O => sig000004cc
    );
  blk00000683 : XORCY
    port map (
      CI => sig000004ce,
      LI => sig000004cd,
      O => sig00000631
    );
  blk00000684 : LUT2
    generic map(
      INIT => X"6"
    )
    port map (
      I0 => sig00000586,
      I1 => sig000006d0,
      O => sig000004cd
    );
  blk00000685 : XORCY
    port map (
      CI => sig000004d0,
      LI => sig000004cf,
      O => sig00000630
    );
  blk00000686 : MUXCY
    port map (
      CI => sig000004d0,
      DI => sig00000586,
      S => sig000004cf,
      O => sig000004ce
    );
  blk00000687 : LUT2
    generic map(
      INIT => X"6"
    )
    port map (
      I0 => sig00000586,
      I1 => sig000006d0,
      O => sig000004cf
    );
  blk00000688 : XORCY
    port map (
      CI => sig000004d2,
      LI => sig000004d1,
      O => sig0000062f
    );
  blk00000689 : MUXCY
    port map (
      CI => sig000004d2,
      DI => sig00000592,
      S => sig000004d1,
      O => sig000004d0
    );
  blk0000068a : LUT2
    generic map(
      INIT => X"6"
    )
    port map (
      I0 => sig00000592,
      I1 => sig000006cf,
      O => sig000004d1
    );
  blk0000068b : XORCY
    port map (
      CI => sig000004d4,
      LI => sig000004d3,
      O => sig0000062e
    );
  blk0000068c : MUXCY
    port map (
      CI => sig000004d4,
      DI => sig00000593,
      S => sig000004d3,
      O => sig000004d2
    );
  blk0000068d : LUT2
    generic map(
      INIT => X"6"
    )
    port map (
      I0 => sig00000593,
      I1 => sig000006ce,
      O => sig000004d3
    );
  blk0000068e : XORCY
    port map (
      CI => sig000004d6,
      LI => sig000004d5,
      O => sig0000062d
    );
  blk0000068f : MUXCY
    port map (
      CI => sig000004d6,
      DI => sig00000594,
      S => sig000004d5,
      O => sig000004d4
    );
  blk00000690 : LUT2
    generic map(
      INIT => X"6"
    )
    port map (
      I0 => sig00000594,
      I1 => sig000006cd,
      O => sig000004d5
    );
  blk00000691 : XORCY
    port map (
      CI => sig000004d8,
      LI => sig000004d7,
      O => sig0000062c
    );
  blk00000692 : MUXCY
    port map (
      CI => sig000004d8,
      DI => sig00000595,
      S => sig000004d7,
      O => sig000004d6
    );
  blk00000693 : LUT2
    generic map(
      INIT => X"6"
    )
    port map (
      I0 => sig00000595,
      I1 => sig000006cc,
      O => sig000004d7
    );
  blk00000694 : XORCY
    port map (
      CI => sig000004da,
      LI => sig000004d9,
      O => sig0000062b
    );
  blk00000695 : MUXCY
    port map (
      CI => sig000004da,
      DI => sig00000596,
      S => sig000004d9,
      O => sig000004d8
    );
  blk00000696 : LUT2
    generic map(
      INIT => X"6"
    )
    port map (
      I0 => sig00000596,
      I1 => sig000006cb,
      O => sig000004d9
    );
  blk00000697 : XORCY
    port map (
      CI => sig000004dc,
      LI => sig000004db,
      O => sig0000062a
    );
  blk00000698 : MUXCY
    port map (
      CI => sig000004dc,
      DI => sig00000597,
      S => sig000004db,
      O => sig000004da
    );
  blk00000699 : LUT2
    generic map(
      INIT => X"6"
    )
    port map (
      I0 => sig00000597,
      I1 => sig000006ca,
      O => sig000004db
    );
  blk0000069a : XORCY
    port map (
      CI => sig000004de,
      LI => sig000004dd,
      O => sig00000629
    );
  blk0000069b : MUXCY
    port map (
      CI => sig000004de,
      DI => sig00000598,
      S => sig000004dd,
      O => sig000004dc
    );
  blk0000069c : LUT2
    generic map(
      INIT => X"6"
    )
    port map (
      I0 => sig00000598,
      I1 => sig000006c9,
      O => sig000004dd
    );
  blk0000069d : XORCY
    port map (
      CI => sig000004e0,
      LI => sig000004df,
      O => sig00000628
    );
  blk0000069e : MUXCY
    port map (
      CI => sig000004e0,
      DI => sig00000599,
      S => sig000004df,
      O => sig000004de
    );
  blk0000069f : LUT2
    generic map(
      INIT => X"6"
    )
    port map (
      I0 => sig00000599,
      I1 => sig000006c8,
      O => sig000004df
    );
  blk000006a0 : XORCY
    port map (
      CI => sig000004e2,
      LI => sig000004e1,
      O => sig00000627
    );
  blk000006a1 : MUXCY
    port map (
      CI => sig000004e2,
      DI => sig0000059a,
      S => sig000004e1,
      O => sig000004e0
    );
  blk000006a2 : LUT2
    generic map(
      INIT => X"6"
    )
    port map (
      I0 => sig0000059a,
      I1 => sig000006c7,
      O => sig000004e1
    );
  blk000006a3 : XORCY
    port map (
      CI => sig000004e4,
      LI => sig000004e3,
      O => sig00000626
    );
  blk000006a4 : MUXCY
    port map (
      CI => sig000004e4,
      DI => sig0000059b,
      S => sig000004e3,
      O => sig000004e2
    );
  blk000006a5 : LUT2
    generic map(
      INIT => X"6"
    )
    port map (
      I0 => sig0000059b,
      I1 => sig000006c6,
      O => sig000004e3
    );
  blk000006a6 : XORCY
    port map (
      CI => sig000004e6,
      LI => sig000004e5,
      O => sig00000625
    );
  blk000006a7 : MUXCY
    port map (
      CI => sig000004e6,
      DI => sig0000059c,
      S => sig000004e5,
      O => sig000004e4
    );
  blk000006a8 : LUT2
    generic map(
      INIT => X"6"
    )
    port map (
      I0 => sig0000059c,
      I1 => sig000006c5,
      O => sig000004e5
    );
  blk000006a9 : XORCY
    port map (
      CI => sig000004e8,
      LI => sig000004e7,
      O => sig00000624
    );
  blk000006aa : MUXCY
    port map (
      CI => sig000004e8,
      DI => sig0000059d,
      S => sig000004e7,
      O => sig000004e6
    );
  blk000006ab : LUT2
    generic map(
      INIT => X"6"
    )
    port map (
      I0 => sig0000059d,
      I1 => sig000006c4,
      O => sig000004e7
    );
  blk000006ac : XORCY
    port map (
      CI => sig000008b6,
      LI => sig000004e9,
      O => sig00000623
    );
  blk000006ad : MUXCY
    port map (
      CI => sig000008b6,
      DI => sig0000059e,
      S => sig000004e9,
      O => sig000004e8
    );
  blk000006ae : LUT2
    generic map(
      INIT => X"6"
    )
    port map (
      I0 => sig0000059e,
      I1 => sig000006c3,
      O => sig000004e9
    );
  blk000006af : XORCY
    port map (
      CI => sig000004eb,
      LI => sig000004ea,
      O => sig00000614
    );
  blk000006b0 : LUT2
    generic map(
      INIT => X"6"
    )
    port map (
      I0 => sig000006c2,
      I1 => sig000006b5,
      O => sig000004ea
    );
  blk000006b1 : XORCY
    port map (
      CI => sig000004ed,
      LI => sig000004ec,
      O => sig00000613
    );
  blk000006b2 : MUXCY
    port map (
      CI => sig000004ed,
      DI => sig000006c2,
      S => sig000004ec,
      O => sig000004eb
    );
  blk000006b3 : LUT2
    generic map(
      INIT => X"6"
    )
    port map (
      I0 => sig000006c2,
      I1 => sig000006b5,
      O => sig000004ec
    );
  blk000006b4 : XORCY
    port map (
      CI => sig000004ef,
      LI => sig000004ee,
      O => sig00000612
    );
  blk000006b5 : MUXCY
    port map (
      CI => sig000004ef,
      DI => sig000006c1,
      S => sig000004ee,
      O => sig000004ed
    );
  blk000006b6 : LUT2
    generic map(
      INIT => X"6"
    )
    port map (
      I0 => sig000006c1,
      I1 => sig000006b4,
      O => sig000004ee
    );
  blk000006b7 : XORCY
    port map (
      CI => sig000004f1,
      LI => sig000004f0,
      O => sig00000611
    );
  blk000006b8 : MUXCY
    port map (
      CI => sig000004f1,
      DI => sig000006c0,
      S => sig000004f0,
      O => sig000004ef
    );
  blk000006b9 : LUT2
    generic map(
      INIT => X"6"
    )
    port map (
      I0 => sig000006c0,
      I1 => sig000006b3,
      O => sig000004f0
    );
  blk000006ba : XORCY
    port map (
      CI => sig000004f3,
      LI => sig000004f2,
      O => sig00000610
    );
  blk000006bb : MUXCY
    port map (
      CI => sig000004f3,
      DI => sig000006bf,
      S => sig000004f2,
      O => sig000004f1
    );
  blk000006bc : LUT2
    generic map(
      INIT => X"6"
    )
    port map (
      I0 => sig000006bf,
      I1 => sig000006b2,
      O => sig000004f2
    );
  blk000006bd : XORCY
    port map (
      CI => sig000004f5,
      LI => sig000004f4,
      O => sig0000060f
    );
  blk000006be : MUXCY
    port map (
      CI => sig000004f5,
      DI => sig000006be,
      S => sig000004f4,
      O => sig000004f3
    );
  blk000006bf : LUT2
    generic map(
      INIT => X"6"
    )
    port map (
      I0 => sig000006be,
      I1 => sig000006b1,
      O => sig000004f4
    );
  blk000006c0 : XORCY
    port map (
      CI => sig000004f7,
      LI => sig000004f6,
      O => sig0000060e
    );
  blk000006c1 : MUXCY
    port map (
      CI => sig000004f7,
      DI => sig000006bd,
      S => sig000004f6,
      O => sig000004f5
    );
  blk000006c2 : LUT2
    generic map(
      INIT => X"6"
    )
    port map (
      I0 => sig000006bd,
      I1 => sig000006b0,
      O => sig000004f6
    );
  blk000006c3 : XORCY
    port map (
      CI => sig000004f9,
      LI => sig000004f8,
      O => sig0000060d
    );
  blk000006c4 : MUXCY
    port map (
      CI => sig000004f9,
      DI => sig000006bc,
      S => sig000004f8,
      O => sig000004f7
    );
  blk000006c5 : LUT2
    generic map(
      INIT => X"6"
    )
    port map (
      I0 => sig000006bc,
      I1 => sig000006af,
      O => sig000004f8
    );
  blk000006c6 : XORCY
    port map (
      CI => sig000004fb,
      LI => sig000004fa,
      O => sig0000060c
    );
  blk000006c7 : MUXCY
    port map (
      CI => sig000004fb,
      DI => sig000006bb,
      S => sig000004fa,
      O => sig000004f9
    );
  blk000006c8 : LUT2
    generic map(
      INIT => X"6"
    )
    port map (
      I0 => sig000006bb,
      I1 => sig000006ae,
      O => sig000004fa
    );
  blk000006c9 : XORCY
    port map (
      CI => sig000004fd,
      LI => sig000004fc,
      O => sig0000060b
    );
  blk000006ca : MUXCY
    port map (
      CI => sig000004fd,
      DI => sig000006ba,
      S => sig000004fc,
      O => sig000004fb
    );
  blk000006cb : LUT2
    generic map(
      INIT => X"6"
    )
    port map (
      I0 => sig000006ba,
      I1 => sig000006ad,
      O => sig000004fc
    );
  blk000006cc : XORCY
    port map (
      CI => sig000004ff,
      LI => sig000004fe,
      O => sig0000060a
    );
  blk000006cd : MUXCY
    port map (
      CI => sig000004ff,
      DI => sig000006b9,
      S => sig000004fe,
      O => sig000004fd
    );
  blk000006ce : LUT2
    generic map(
      INIT => X"6"
    )
    port map (
      I0 => sig000006b9,
      I1 => sig000006ac,
      O => sig000004fe
    );
  blk000006cf : XORCY
    port map (
      CI => sig00000501,
      LI => sig00000500,
      O => sig00000609
    );
  blk000006d0 : MUXCY
    port map (
      CI => sig00000501,
      DI => sig000006b8,
      S => sig00000500,
      O => sig000004ff
    );
  blk000006d1 : LUT2
    generic map(
      INIT => X"6"
    )
    port map (
      I0 => sig000006b8,
      I1 => sig000006ab,
      O => sig00000500
    );
  blk000006d2 : XORCY
    port map (
      CI => sig00000503,
      LI => sig00000502,
      O => sig00000608
    );
  blk000006d3 : MUXCY
    port map (
      CI => sig00000503,
      DI => sig000006b7,
      S => sig00000502,
      O => sig00000501
    );
  blk000006d4 : LUT2
    generic map(
      INIT => X"6"
    )
    port map (
      I0 => sig000006b7,
      I1 => sig000006aa,
      O => sig00000502
    );
  blk000006d5 : XORCY
    port map (
      CI => sig000008b6,
      LI => sig00000504,
      O => sig00000607
    );
  blk000006d6 : MUXCY
    port map (
      CI => sig000008b6,
      DI => sig000006b6,
      S => sig00000504,
      O => sig00000503
    );
  blk000006d7 : LUT2
    generic map(
      INIT => X"6"
    )
    port map (
      I0 => sig000006b6,
      I1 => sig000006a9,
      O => sig00000504
    );
  blk000006d8 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => sig00000631,
      Q => sig00000635
    );
  blk000006d9 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => sig00000630,
      Q => sig00000634
    );
  blk000006da : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => sig0000062f,
      Q => sig00000633
    );
  blk000006db : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => sig0000062e,
      Q => sig00000632
    );
  blk000006dc : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => sig00000622,
      Q => sig00000639
    );
  blk000006dd : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => sig00000621,
      Q => sig00000638
    );
  blk000006de : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => sig00000620,
      Q => sig00000637
    );
  blk000006df : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => sig0000061f,
      Q => sig00000636
    );
  blk000006e0 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => sig00000614,
      Q => sig0000059f
    );
  blk000006e1 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => sig00000613,
      Q => sig000005a4
    );
  blk000006e2 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => sig00000612,
      Q => sig000005a5
    );
  blk000006e3 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => sig00000611,
      Q => sig000005a6
    );
  blk000006e4 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => sig00000610,
      Q => sig000005a7
    );
  blk000006e5 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => sig0000060f,
      Q => sig000005a8
    );
  blk000006e6 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => sig0000060e,
      Q => sig000005a9
    );
  blk000006e7 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => sig0000060d,
      Q => sig000005aa
    );
  blk000006e8 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => sig0000060c,
      Q => sig000005ab
    );
  blk000006e9 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => sig0000060b,
      Q => sig000005ac
    );
  blk000006ea : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => sig0000060a,
      Q => sig000005ad
    );
  blk000006eb : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => sig00000609,
      Q => sig000005ae
    );
  blk000006ec : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => sig00000608,
      Q => sig000005af
    );
  blk000006ed : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => sig00000607,
      Q => sig000005b0
    );
  blk000006ee : XORCY
    port map (
      CI => sig000006d2,
      LI => sig000006d1,
      O => sig0000071b
    );
  blk000006ef : XORCY
    port map (
      CI => sig000006d4,
      LI => sig000006d3,
      O => sig0000071a
    );
  blk000006f0 : MUXCY
    port map (
      CI => sig000006d4,
      DI => sig000008b6,
      S => sig000006d3,
      O => sig000006d2
    );
  blk000006f1 : XORCY
    port map (
      CI => sig000006d6,
      LI => sig000006d5,
      O => sig00000719
    );
  blk000006f2 : MUXCY
    port map (
      CI => sig000006d6,
      DI => sig000008b6,
      S => sig000006d5,
      O => sig000006d4
    );
  blk000006f3 : XORCY
    port map (
      CI => sig000006d8,
      LI => sig000006d7,
      O => sig00000718
    );
  blk000006f4 : MUXCY
    port map (
      CI => sig000006d8,
      DI => sig000008b6,
      S => sig000006d7,
      O => sig000006d6
    );
  blk000006f5 : XORCY
    port map (
      CI => sig000006da,
      LI => sig000006d9,
      O => sig00000717
    );
  blk000006f6 : MUXCY
    port map (
      CI => sig000006da,
      DI => sig000008b6,
      S => sig000006d9,
      O => sig000006d8
    );
  blk000006f7 : XORCY
    port map (
      CI => sig000006dc,
      LI => sig000006db,
      O => sig00000716
    );
  blk000006f8 : MUXCY
    port map (
      CI => sig000006dc,
      DI => sig000008b6,
      S => sig000006db,
      O => sig000006da
    );
  blk000006f9 : XORCY
    port map (
      CI => sig000006de,
      LI => sig000006dd,
      O => sig00000715
    );
  blk000006fa : MUXCY
    port map (
      CI => sig000006de,
      DI => sig000008b6,
      S => sig000006dd,
      O => sig000006dc
    );
  blk000006fb : XORCY
    port map (
      CI => sig000006e0,
      LI => sig000006df,
      O => sig00000714
    );
  blk000006fc : MUXCY
    port map (
      CI => sig000006e0,
      DI => sig000008b6,
      S => sig000006df,
      O => sig000006de
    );
  blk000006fd : XORCY
    port map (
      CI => sig000006e2,
      LI => sig000006e1,
      O => sig00000713
    );
  blk000006fe : MUXCY
    port map (
      CI => sig000006e2,
      DI => sig000008b6,
      S => sig000006e1,
      O => sig000006e0
    );
  blk000006ff : XORCY
    port map (
      CI => sig000006e4,
      LI => sig000006e3,
      O => sig00000712
    );
  blk00000700 : MUXCY
    port map (
      CI => sig000006e4,
      DI => sig000008b6,
      S => sig000006e3,
      O => sig000006e2
    );
  blk00000701 : XORCY
    port map (
      CI => sig000006e6,
      LI => sig000006e5,
      O => sig00000711
    );
  blk00000702 : MUXCY
    port map (
      CI => sig000006e6,
      DI => sig000008b6,
      S => sig000006e5,
      O => sig000006e4
    );
  blk00000703 : XORCY
    port map (
      CI => sig000006e8,
      LI => sig000006e7,
      O => sig00000710
    );
  blk00000704 : MUXCY
    port map (
      CI => sig000006e8,
      DI => sig000008b6,
      S => sig000006e7,
      O => sig000006e6
    );
  blk00000705 : XORCY
    port map (
      CI => sig000006d1,
      LI => sig000006e9,
      O => sig0000070f
    );
  blk00000706 : MUXCY
    port map (
      CI => sig000006d1,
      DI => sig000008b6,
      S => sig000006e9,
      O => sig000006e8
    );
  blk00000707 : XORCY
    port map (
      CI => sig000006ea,
      LI => sig000006d1,
      O => sig00000735
    );
  blk00000708 : XORCY
    port map (
      CI => sig000006ec,
      LI => sig000006eb,
      O => sig00000734
    );
  blk00000709 : MUXCY
    port map (
      CI => sig000006ec,
      DI => sig000008b6,
      S => sig000006eb,
      O => sig000006ea
    );
  blk0000070a : XORCY
    port map (
      CI => sig000006ee,
      LI => sig000006ed,
      O => sig00000733
    );
  blk0000070b : MUXCY
    port map (
      CI => sig000006ee,
      DI => sig000008b6,
      S => sig000006ed,
      O => sig000006ec
    );
  blk0000070c : XORCY
    port map (
      CI => sig000006f0,
      LI => sig000006ef,
      O => sig00000732
    );
  blk0000070d : MUXCY
    port map (
      CI => sig000006f0,
      DI => sig000008b6,
      S => sig000006ef,
      O => sig000006ee
    );
  blk0000070e : XORCY
    port map (
      CI => sig000006f2,
      LI => sig000006f1,
      O => sig00000731
    );
  blk0000070f : MUXCY
    port map (
      CI => sig000006f2,
      DI => sig000008b6,
      S => sig000006f1,
      O => sig000006f0
    );
  blk00000710 : XORCY
    port map (
      CI => sig000006f4,
      LI => sig000006f3,
      O => sig00000730
    );
  blk00000711 : MUXCY
    port map (
      CI => sig000006f4,
      DI => sig000008b6,
      S => sig000006f3,
      O => sig000006f2
    );
  blk00000712 : XORCY
    port map (
      CI => sig000006f6,
      LI => sig000006f5,
      O => sig0000072f
    );
  blk00000713 : MUXCY
    port map (
      CI => sig000006f6,
      DI => sig000008b6,
      S => sig000006f5,
      O => sig000006f4
    );
  blk00000714 : XORCY
    port map (
      CI => sig000006f8,
      LI => sig000006f7,
      O => sig0000072e
    );
  blk00000715 : MUXCY
    port map (
      CI => sig000006f8,
      DI => sig000008b6,
      S => sig000006f7,
      O => sig000006f6
    );
  blk00000716 : XORCY
    port map (
      CI => sig000006fa,
      LI => sig000006f9,
      O => sig0000072d
    );
  blk00000717 : MUXCY
    port map (
      CI => sig000006fa,
      DI => sig000008b6,
      S => sig000006f9,
      O => sig000006f8
    );
  blk00000718 : XORCY
    port map (
      CI => sig000006fc,
      LI => sig000006fb,
      O => sig0000072c
    );
  blk00000719 : MUXCY
    port map (
      CI => sig000006fc,
      DI => sig000008b6,
      S => sig000006fb,
      O => sig000006fa
    );
  blk0000071a : XORCY
    port map (
      CI => sig000006fe,
      LI => sig000006fd,
      O => sig0000072b
    );
  blk0000071b : MUXCY
    port map (
      CI => sig000006fe,
      DI => sig000008b6,
      S => sig000006fd,
      O => sig000006fc
    );
  blk0000071c : XORCY
    port map (
      CI => sig00000700,
      LI => sig000006ff,
      O => sig0000072a
    );
  blk0000071d : MUXCY
    port map (
      CI => sig00000700,
      DI => sig000008b6,
      S => sig000006ff,
      O => sig000006fe
    );
  blk0000071e : XORCY
    port map (
      CI => sig000006d1,
      LI => sig00000701,
      O => sig00000729
    );
  blk0000071f : MUXCY
    port map (
      CI => sig000006d1,
      DI => sig000008b6,
      S => sig00000701,
      O => sig00000700
    );
  blk00000720 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => sig00000728,
      Q => sig000006c2
    );
  blk00000721 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => sig00000727,
      Q => sig000006c1
    );
  blk00000722 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => sig00000726,
      Q => sig000006c0
    );
  blk00000723 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => sig00000725,
      Q => sig000006bf
    );
  blk00000724 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => sig00000724,
      Q => sig000006be
    );
  blk00000725 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => sig00000723,
      Q => sig000006bd
    );
  blk00000726 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => sig00000722,
      Q => sig000006bc
    );
  blk00000727 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => sig00000721,
      Q => sig000006bb
    );
  blk00000728 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => sig00000720,
      Q => sig000006ba
    );
  blk00000729 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => sig0000071f,
      Q => sig000006b9
    );
  blk0000072a : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => sig0000071e,
      Q => sig000006b8
    );
  blk0000072b : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => sig0000071d,
      Q => sig000006b7
    );
  blk0000072c : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => sig0000071c,
      Q => sig000006b6
    );
  blk0000072d : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => sig0000070e,
      Q => sig000006b5
    );
  blk0000072e : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => sig0000070d,
      Q => sig000006b4
    );
  blk0000072f : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => sig0000070c,
      Q => sig000006b3
    );
  blk00000730 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => sig0000070b,
      Q => sig000006b2
    );
  blk00000731 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => sig0000070a,
      Q => sig000006b1
    );
  blk00000732 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => sig00000709,
      Q => sig000006b0
    );
  blk00000733 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => sig00000708,
      Q => sig000006af
    );
  blk00000734 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => sig00000707,
      Q => sig000006ae
    );
  blk00000735 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => sig00000706,
      Q => sig000006ad
    );
  blk00000736 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => sig00000705,
      Q => sig000006ac
    );
  blk00000737 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => sig00000704,
      Q => sig000006ab
    );
  blk00000738 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => sig00000703,
      Q => sig000006aa
    );
  blk00000739 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => sig00000702,
      Q => sig000006a9
    );
  blk0000073a : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => sig00000240,
      Q => sig000006d0
    );
  blk0000073b : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => sig0000023f,
      Q => sig000006cf
    );
  blk0000073c : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => sig0000023e,
      Q => sig000006ce
    );
  blk0000073d : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => sig0000023d,
      Q => sig000006cd
    );
  blk0000073e : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => sig0000023c,
      Q => sig000006cc
    );
  blk0000073f : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => sig0000023b,
      Q => sig000006cb
    );
  blk00000740 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => sig0000023a,
      Q => sig000006ca
    );
  blk00000741 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => sig00000239,
      Q => sig000006c9
    );
  blk00000742 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => sig00000238,
      Q => sig000006c8
    );
  blk00000743 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => sig00000237,
      Q => sig000006c7
    );
  blk00000744 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => sig00000236,
      Q => sig000006c6
    );
  blk00000745 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => sig00000235,
      Q => sig000006c5
    );
  blk00000746 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => sig00000234,
      Q => sig000006c4
    );
  blk00000747 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => sig00000233,
      Q => sig000006c3
    );
  blk00000748 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => sig0000024e,
      Q => sig00000586
    );
  blk00000749 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => sig0000024d,
      Q => sig00000592
    );
  blk0000074a : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => sig0000024c,
      Q => sig00000593
    );
  blk0000074b : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => sig0000024b,
      Q => sig00000594
    );
  blk0000074c : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => sig0000024a,
      Q => sig00000595
    );
  blk0000074d : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => sig00000249,
      Q => sig00000596
    );
  blk0000074e : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => sig00000248,
      Q => sig00000597
    );
  blk0000074f : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => sig00000247,
      Q => sig00000598
    );
  blk00000750 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => sig00000246,
      Q => sig00000599
    );
  blk00000751 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => sig00000245,
      Q => sig0000059a
    );
  blk00000752 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => sig00000244,
      Q => sig0000059b
    );
  blk00000753 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => sig00000243,
      Q => sig0000059c
    );
  blk00000754 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => sig00000242,
      Q => sig0000059d
    );
  blk00000755 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => sig00000241,
      Q => sig0000059e
    );
  blk00000756 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => sig00000639,
      Q => sig00000549
    );
  blk00000757 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => sig00000638,
      Q => sig0000054d
    );
  blk00000758 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => sig00000637,
      Q => sig0000054e
    );
  blk00000759 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => sig00000636,
      Q => sig0000054f
    );
  blk0000075a : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => sig00000635,
      Q => sig000005f5
    );
  blk0000075b : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => sig00000634,
      Q => sig000005f9
    );
  blk0000075c : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => sig00000633,
      Q => sig000005fa
    );
  blk0000075d : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => sig00000632,
      Q => sig000005fb
    );
  blk00000767 : LUT6
    generic map(
      INIT => X"FF00F0F0CCCCAAAA"
    )
    port map (
      I0 => sig000008b6,
      I1 => sig000008b6,
      I2 => sig000008b6,
      I3 => sig00000200,
      I4 => sig00000251,
      I5 => sig00000252,
      O => sig00000736
    );
  blk00000768 : LUT6
    generic map(
      INIT => X"FF00F0F0CCCCAAAA"
    )
    port map (
      I0 => sig000008b6,
      I1 => sig000008b6,
      I2 => sig00000200,
      I3 => sig00000201,
      I4 => sig00000251,
      I5 => sig00000252,
      O => sig00000737
    );
  blk00000769 : LUT6
    generic map(
      INIT => X"FF00F0F0CCCCAAAA"
    )
    port map (
      I0 => sig000008b6,
      I1 => sig00000200,
      I2 => sig00000201,
      I3 => sig00000202,
      I4 => sig00000251,
      I5 => sig00000252,
      O => sig00000738
    );
  blk0000076a : LUT6
    generic map(
      INIT => X"FF00F0F0CCCCAAAA"
    )
    port map (
      I0 => sig00000200,
      I1 => sig00000201,
      I2 => sig00000202,
      I3 => sig00000203,
      I4 => sig00000251,
      I5 => sig00000252,
      O => sig00000739
    );
  blk0000076b : LUT6
    generic map(
      INIT => X"FF00F0F0CCCCAAAA"
    )
    port map (
      I0 => sig00000201,
      I1 => sig00000202,
      I2 => sig00000203,
      I3 => sig00000204,
      I4 => sig00000251,
      I5 => sig00000252,
      O => sig0000073a
    );
  blk0000076c : LUT6
    generic map(
      INIT => X"FF00F0F0CCCCAAAA"
    )
    port map (
      I0 => sig00000202,
      I1 => sig00000203,
      I2 => sig00000204,
      I3 => sig00000205,
      I4 => sig00000251,
      I5 => sig00000252,
      O => sig0000073b
    );
  blk0000076d : LUT6
    generic map(
      INIT => X"FF00F0F0CCCCAAAA"
    )
    port map (
      I0 => sig00000203,
      I1 => sig00000204,
      I2 => sig00000205,
      I3 => sig00000206,
      I4 => sig00000251,
      I5 => sig00000252,
      O => sig0000073c
    );
  blk0000076e : LUT6
    generic map(
      INIT => X"FF00F0F0CCCCAAAA"
    )
    port map (
      I0 => sig00000204,
      I1 => sig00000205,
      I2 => sig00000206,
      I3 => sig00000207,
      I4 => sig00000251,
      I5 => sig00000252,
      O => sig0000073d
    );
  blk0000076f : LUT6
    generic map(
      INIT => X"FF00F0F0CCCCAAAA"
    )
    port map (
      I0 => sig00000205,
      I1 => sig00000206,
      I2 => sig00000207,
      I3 => sig00000208,
      I4 => sig00000251,
      I5 => sig00000252,
      O => sig0000073e
    );
  blk00000770 : LUT6
    generic map(
      INIT => X"FF00F0F0CCCCAAAA"
    )
    port map (
      I0 => sig00000206,
      I1 => sig00000207,
      I2 => sig00000208,
      I3 => sig00000209,
      I4 => sig00000251,
      I5 => sig00000252,
      O => sig0000073f
    );
  blk00000771 : LUT6
    generic map(
      INIT => X"FF00F0F0CCCCAAAA"
    )
    port map (
      I0 => sig00000207,
      I1 => sig00000208,
      I2 => sig00000209,
      I3 => sig0000020a,
      I4 => sig00000251,
      I5 => sig00000252,
      O => sig00000740
    );
  blk00000772 : LUT6
    generic map(
      INIT => X"FF00F0F0CCCCAAAA"
    )
    port map (
      I0 => sig00000208,
      I1 => sig00000209,
      I2 => sig0000020a,
      I3 => sig0000020b,
      I4 => sig00000251,
      I5 => sig00000252,
      O => sig00000741
    );
  blk00000773 : LUT6
    generic map(
      INIT => X"FF00F0F0CCCCAAAA"
    )
    port map (
      I0 => sig00000209,
      I1 => sig0000020a,
      I2 => sig0000020b,
      I3 => sig0000020c,
      I4 => sig00000251,
      I5 => sig00000252,
      O => sig00000742
    );
  blk00000774 : LUT6
    generic map(
      INIT => X"FF00F0F0CCCCAAAA"
    )
    port map (
      I0 => sig0000020a,
      I1 => sig0000020b,
      I2 => sig0000020c,
      I3 => sig0000020d,
      I4 => sig00000251,
      I5 => sig00000252,
      O => sig00000743
    );
  blk00000775 : LUT6
    generic map(
      INIT => X"FF00F0F0CCCCAAAA"
    )
    port map (
      I0 => sig0000020b,
      I1 => sig0000020c,
      I2 => sig0000020d,
      I3 => sig0000020e,
      I4 => sig00000251,
      I5 => sig00000252,
      O => sig00000744
    );
  blk00000776 : LUT6
    generic map(
      INIT => X"FF00F0F0CCCCAAAA"
    )
    port map (
      I0 => sig0000020c,
      I1 => sig0000020d,
      I2 => sig0000020e,
      I3 => sig0000020f,
      I4 => sig00000251,
      I5 => sig00000252,
      O => sig00000745
    );
  blk00000777 : LUT6
    generic map(
      INIT => X"FF00F0F0CCCCAAAA"
    )
    port map (
      I0 => sig0000020d,
      I1 => sig0000020e,
      I2 => sig0000020f,
      I3 => sig00000210,
      I4 => sig00000251,
      I5 => sig00000252,
      O => sig00000746
    );
  blk00000778 : LUT6
    generic map(
      INIT => X"FF00F0F0CCCCAAAA"
    )
    port map (
      I0 => sig0000020e,
      I1 => sig0000020f,
      I2 => sig00000210,
      I3 => sig00000211,
      I4 => sig00000251,
      I5 => sig00000252,
      O => sig00000747
    );
  blk00000779 : LUT6
    generic map(
      INIT => X"FF00F0F0CCCCAAAA"
    )
    port map (
      I0 => sig0000020f,
      I1 => sig00000210,
      I2 => sig00000211,
      I3 => sig00000212,
      I4 => sig00000251,
      I5 => sig00000252,
      O => sig00000748
    );
  blk0000077a : LUT6
    generic map(
      INIT => X"FF00F0F0CCCCAAAA"
    )
    port map (
      I0 => sig00000210,
      I1 => sig00000211,
      I2 => sig00000212,
      I3 => sig00000213,
      I4 => sig00000251,
      I5 => sig00000252,
      O => sig00000749
    );
  blk0000077b : LUT6
    generic map(
      INIT => X"FF00F0F0CCCCAAAA"
    )
    port map (
      I0 => sig00000211,
      I1 => sig00000212,
      I2 => sig00000213,
      I3 => sig00000213,
      I4 => sig00000251,
      I5 => sig00000252,
      O => sig0000074a
    );
  blk0000077c : LUT6
    generic map(
      INIT => X"FF00F0F0CCCCAAAA"
    )
    port map (
      I0 => sig00000212,
      I1 => sig00000213,
      I2 => sig00000213,
      I3 => sig00000213,
      I4 => sig00000251,
      I5 => sig00000252,
      O => sig0000074b
    );
  blk0000077d : LUT6
    generic map(
      INIT => X"FF00F0F0CCCCAAAA"
    )
    port map (
      I0 => sig00000213,
      I1 => sig00000213,
      I2 => sig00000213,
      I3 => sig00000213,
      I4 => sig00000251,
      I5 => sig00000252,
      O => sig0000074c
    );
  blk0000077e : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => sig00000736,
      R => sig000008b6,
      Q => NLW_blk0000077e_Q_UNCONNECTED
    );
  blk0000077f : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => sig00000737,
      R => sig000008b6,
      Q => NLW_blk0000077f_Q_UNCONNECTED
    );
  blk00000780 : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => sig00000738,
      R => sig000008b6,
      Q => NLW_blk00000780_Q_UNCONNECTED
    );
  blk00000781 : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => sig00000739,
      R => sig000008b6,
      Q => NLW_blk00000781_Q_UNCONNECTED
    );
  blk00000782 : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => sig0000073a,
      R => sig000008b6,
      Q => NLW_blk00000782_Q_UNCONNECTED
    );
  blk00000783 : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => sig0000073b,
      R => sig000008b6,
      Q => NLW_blk00000783_Q_UNCONNECTED
    );
  blk00000784 : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => sig0000073c,
      R => sig000008b6,
      Q => NLW_blk00000784_Q_UNCONNECTED
    );
  blk00000785 : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => sig0000073d,
      R => sig000008b6,
      Q => NLW_blk00000785_Q_UNCONNECTED
    );
  blk00000786 : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => sig0000073e,
      R => sig000008b6,
      Q => sig000000fb
    );
  blk00000787 : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => sig0000073f,
      R => sig000008b6,
      Q => sig000000fc
    );
  blk00000788 : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => sig00000740,
      R => sig000008b6,
      Q => sig000000fd
    );
  blk00000789 : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => sig00000741,
      R => sig000008b6,
      Q => sig000000fe
    );
  blk0000078a : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => sig00000742,
      R => sig000008b6,
      Q => sig000000ff
    );
  blk0000078b : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => sig00000743,
      R => sig000008b6,
      Q => sig00000100
    );
  blk0000078c : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => sig00000744,
      R => sig000008b6,
      Q => sig00000101
    );
  blk0000078d : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => sig00000745,
      R => sig000008b6,
      Q => sig00000102
    );
  blk0000078e : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => sig00000746,
      R => sig000008b6,
      Q => sig00000103
    );
  blk0000078f : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => sig00000747,
      R => sig000008b6,
      Q => sig00000104
    );
  blk00000790 : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => sig00000748,
      R => sig000008b6,
      Q => sig00000105
    );
  blk00000791 : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => sig00000749,
      R => sig000008b6,
      Q => sig00000106
    );
  blk00000792 : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => sig0000074a,
      R => sig000008b6,
      Q => NLW_blk00000792_Q_UNCONNECTED
    );
  blk00000793 : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => sig0000074b,
      R => sig000008b6,
      Q => NLW_blk00000793_Q_UNCONNECTED
    );
  blk00000794 : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => sig0000074c,
      R => sig000008b6,
      Q => NLW_blk00000794_Q_UNCONNECTED
    );
  blk00000795 : LUT6
    generic map(
      INIT => X"FF00F0F0CCCCAAAA"
    )
    port map (
      I0 => sig000008b6,
      I1 => sig000008b6,
      I2 => sig000008b6,
      I3 => sig000001ec,
      I4 => sig00000251,
      I5 => sig00000252,
      O => sig0000074d
    );
  blk00000796 : LUT6
    generic map(
      INIT => X"FF00F0F0CCCCAAAA"
    )
    port map (
      I0 => sig000008b6,
      I1 => sig000008b6,
      I2 => sig000001ec,
      I3 => sig000001ed,
      I4 => sig00000251,
      I5 => sig00000252,
      O => sig0000074e
    );
  blk00000797 : LUT6
    generic map(
      INIT => X"FF00F0F0CCCCAAAA"
    )
    port map (
      I0 => sig000008b6,
      I1 => sig000001ec,
      I2 => sig000001ed,
      I3 => sig000001ee,
      I4 => sig00000251,
      I5 => sig00000252,
      O => sig0000074f
    );
  blk00000798 : LUT6
    generic map(
      INIT => X"FF00F0F0CCCCAAAA"
    )
    port map (
      I0 => sig000001ec,
      I1 => sig000001ed,
      I2 => sig000001ee,
      I3 => sig000001ef,
      I4 => sig00000251,
      I5 => sig00000252,
      O => sig00000750
    );
  blk00000799 : LUT6
    generic map(
      INIT => X"FF00F0F0CCCCAAAA"
    )
    port map (
      I0 => sig000001ed,
      I1 => sig000001ee,
      I2 => sig000001ef,
      I3 => sig000001f0,
      I4 => sig00000251,
      I5 => sig00000252,
      O => sig00000751
    );
  blk0000079a : LUT6
    generic map(
      INIT => X"FF00F0F0CCCCAAAA"
    )
    port map (
      I0 => sig000001ee,
      I1 => sig000001ef,
      I2 => sig000001f0,
      I3 => sig000001f1,
      I4 => sig00000251,
      I5 => sig00000252,
      O => sig00000752
    );
  blk0000079b : LUT6
    generic map(
      INIT => X"FF00F0F0CCCCAAAA"
    )
    port map (
      I0 => sig000001ef,
      I1 => sig000001f0,
      I2 => sig000001f1,
      I3 => sig000001f2,
      I4 => sig00000251,
      I5 => sig00000252,
      O => sig00000753
    );
  blk0000079c : LUT6
    generic map(
      INIT => X"FF00F0F0CCCCAAAA"
    )
    port map (
      I0 => sig000001f0,
      I1 => sig000001f1,
      I2 => sig000001f2,
      I3 => sig000001f3,
      I4 => sig00000251,
      I5 => sig00000252,
      O => sig00000754
    );
  blk0000079d : LUT6
    generic map(
      INIT => X"FF00F0F0CCCCAAAA"
    )
    port map (
      I0 => sig000001f1,
      I1 => sig000001f2,
      I2 => sig000001f3,
      I3 => sig000001f4,
      I4 => sig00000251,
      I5 => sig00000252,
      O => sig00000755
    );
  blk0000079e : LUT6
    generic map(
      INIT => X"FF00F0F0CCCCAAAA"
    )
    port map (
      I0 => sig000001f2,
      I1 => sig000001f3,
      I2 => sig000001f4,
      I3 => sig000001f5,
      I4 => sig00000251,
      I5 => sig00000252,
      O => sig00000756
    );
  blk0000079f : LUT6
    generic map(
      INIT => X"FF00F0F0CCCCAAAA"
    )
    port map (
      I0 => sig000001f3,
      I1 => sig000001f4,
      I2 => sig000001f5,
      I3 => sig000001f6,
      I4 => sig00000251,
      I5 => sig00000252,
      O => sig00000757
    );
  blk000007a0 : LUT6
    generic map(
      INIT => X"FF00F0F0CCCCAAAA"
    )
    port map (
      I0 => sig000001f4,
      I1 => sig000001f5,
      I2 => sig000001f6,
      I3 => sig000001f7,
      I4 => sig00000251,
      I5 => sig00000252,
      O => sig00000758
    );
  blk000007a1 : LUT6
    generic map(
      INIT => X"FF00F0F0CCCCAAAA"
    )
    port map (
      I0 => sig000001f5,
      I1 => sig000001f6,
      I2 => sig000001f7,
      I3 => sig000001f8,
      I4 => sig00000251,
      I5 => sig00000252,
      O => sig00000759
    );
  blk000007a2 : LUT6
    generic map(
      INIT => X"FF00F0F0CCCCAAAA"
    )
    port map (
      I0 => sig000001f6,
      I1 => sig000001f7,
      I2 => sig000001f8,
      I3 => sig000001f9,
      I4 => sig00000251,
      I5 => sig00000252,
      O => sig0000075a
    );
  blk000007a3 : LUT6
    generic map(
      INIT => X"FF00F0F0CCCCAAAA"
    )
    port map (
      I0 => sig000001f7,
      I1 => sig000001f8,
      I2 => sig000001f9,
      I3 => sig000001fa,
      I4 => sig00000251,
      I5 => sig00000252,
      O => sig0000075b
    );
  blk000007a4 : LUT6
    generic map(
      INIT => X"FF00F0F0CCCCAAAA"
    )
    port map (
      I0 => sig000001f8,
      I1 => sig000001f9,
      I2 => sig000001fa,
      I3 => sig000001fb,
      I4 => sig00000251,
      I5 => sig00000252,
      O => sig0000075c
    );
  blk000007a5 : LUT6
    generic map(
      INIT => X"FF00F0F0CCCCAAAA"
    )
    port map (
      I0 => sig000001f9,
      I1 => sig000001fa,
      I2 => sig000001fb,
      I3 => sig000001fc,
      I4 => sig00000251,
      I5 => sig00000252,
      O => sig0000075d
    );
  blk000007a6 : LUT6
    generic map(
      INIT => X"FF00F0F0CCCCAAAA"
    )
    port map (
      I0 => sig000001fa,
      I1 => sig000001fb,
      I2 => sig000001fc,
      I3 => sig000001fd,
      I4 => sig00000251,
      I5 => sig00000252,
      O => sig0000075e
    );
  blk000007a7 : LUT6
    generic map(
      INIT => X"FF00F0F0CCCCAAAA"
    )
    port map (
      I0 => sig000001fb,
      I1 => sig000001fc,
      I2 => sig000001fd,
      I3 => sig000001fe,
      I4 => sig00000251,
      I5 => sig00000252,
      O => sig0000075f
    );
  blk000007a8 : LUT6
    generic map(
      INIT => X"FF00F0F0CCCCAAAA"
    )
    port map (
      I0 => sig000001fc,
      I1 => sig000001fd,
      I2 => sig000001fe,
      I3 => sig000001ff,
      I4 => sig00000251,
      I5 => sig00000252,
      O => sig00000760
    );
  blk000007a9 : LUT6
    generic map(
      INIT => X"FF00F0F0CCCCAAAA"
    )
    port map (
      I0 => sig000001fd,
      I1 => sig000001fe,
      I2 => sig000001ff,
      I3 => sig000001ff,
      I4 => sig00000251,
      I5 => sig00000252,
      O => sig00000761
    );
  blk000007aa : LUT6
    generic map(
      INIT => X"FF00F0F0CCCCAAAA"
    )
    port map (
      I0 => sig000001fe,
      I1 => sig000001ff,
      I2 => sig000001ff,
      I3 => sig000001ff,
      I4 => sig00000251,
      I5 => sig00000252,
      O => sig00000762
    );
  blk000007ab : LUT6
    generic map(
      INIT => X"FF00F0F0CCCCAAAA"
    )
    port map (
      I0 => sig000001ff,
      I1 => sig000001ff,
      I2 => sig000001ff,
      I3 => sig000001ff,
      I4 => sig00000251,
      I5 => sig00000252,
      O => sig00000763
    );
  blk000007ac : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => sig0000074d,
      R => sig000008b6,
      Q => NLW_blk000007ac_Q_UNCONNECTED
    );
  blk000007ad : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => sig0000074e,
      R => sig000008b6,
      Q => NLW_blk000007ad_Q_UNCONNECTED
    );
  blk000007ae : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => sig0000074f,
      R => sig000008b6,
      Q => NLW_blk000007ae_Q_UNCONNECTED
    );
  blk000007af : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => sig00000750,
      R => sig000008b6,
      Q => NLW_blk000007af_Q_UNCONNECTED
    );
  blk000007b0 : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => sig00000751,
      R => sig000008b6,
      Q => NLW_blk000007b0_Q_UNCONNECTED
    );
  blk000007b1 : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => sig00000752,
      R => sig000008b6,
      Q => NLW_blk000007b1_Q_UNCONNECTED
    );
  blk000007b2 : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => sig00000753,
      R => sig000008b6,
      Q => NLW_blk000007b2_Q_UNCONNECTED
    );
  blk000007b3 : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => sig00000754,
      R => sig000008b6,
      Q => NLW_blk000007b3_Q_UNCONNECTED
    );
  blk000007b4 : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => sig00000755,
      R => sig000008b6,
      Q => sig000000ef
    );
  blk000007b5 : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => sig00000756,
      R => sig000008b6,
      Q => sig000000f0
    );
  blk000007b6 : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => sig00000757,
      R => sig000008b6,
      Q => sig000000f1
    );
  blk000007b7 : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => sig00000758,
      R => sig000008b6,
      Q => sig000000f2
    );
  blk000007b8 : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => sig00000759,
      R => sig000008b6,
      Q => sig000000f3
    );
  blk000007b9 : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => sig0000075a,
      R => sig000008b6,
      Q => sig000000f4
    );
  blk000007ba : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => sig0000075b,
      R => sig000008b6,
      Q => sig000000f5
    );
  blk000007bb : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => sig0000075c,
      R => sig000008b6,
      Q => sig000000f6
    );
  blk000007bc : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => sig0000075d,
      R => sig000008b6,
      Q => sig000000f7
    );
  blk000007bd : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => sig0000075e,
      R => sig000008b6,
      Q => sig000000f8
    );
  blk000007be : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => sig0000075f,
      R => sig000008b6,
      Q => sig000000f9
    );
  blk000007bf : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => sig00000760,
      R => sig000008b6,
      Q => sig000000fa
    );
  blk000007c0 : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => sig00000761,
      R => sig000008b6,
      Q => NLW_blk000007c0_Q_UNCONNECTED
    );
  blk000007c1 : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => sig00000762,
      R => sig000008b6,
      Q => NLW_blk000007c1_Q_UNCONNECTED
    );
  blk000007c2 : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => sig00000763,
      R => sig000008b6,
      Q => NLW_blk000007c2_Q_UNCONNECTED
    );
  blk000007c3 : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => sig00000764,
      R => sig000008b6,
      Q => NLW_blk000007c3_Q_UNCONNECTED
    );
  blk000007c4 : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => sig00000765,
      R => sig000008b6,
      Q => NLW_blk000007c4_Q_UNCONNECTED
    );
  blk000007c5 : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => sig00000766,
      R => sig000008b6,
      Q => NLW_blk000007c5_Q_UNCONNECTED
    );
  blk000007c6 : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => sig00000767,
      R => sig000008b6,
      Q => sig000000d6
    );
  blk000007c7 : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => sig00000768,
      R => sig000008b6,
      Q => sig000000d5
    );
  blk000007c8 : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => sig00000769,
      R => sig000008b6,
      Q => sig000000d4
    );
  blk000007c9 : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => sig0000076a,
      R => sig000008b6,
      Q => sig000000d3
    );
  blk000007ca : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => sig0000076b,
      R => sig000008b6,
      Q => sig000000d2
    );
  blk000007cb : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => sig0000076c,
      R => sig000008b6,
      Q => sig000000d1
    );
  blk000007cc : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => sig0000076d,
      R => sig000008b6,
      Q => sig000000d0
    );
  blk000007cd : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => sig0000076e,
      R => sig000008b6,
      Q => sig000000cf
    );
  blk000007ce : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => sig0000076f,
      R => sig000008b6,
      Q => sig000000ce
    );
  blk000007cf : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => sig00000770,
      R => sig000008b6,
      Q => sig000000cd
    );
  blk000007d0 : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => sig00000771,
      R => sig000008b6,
      Q => sig000000cc
    );
  blk000007d1 : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => sig00000772,
      R => sig000008b6,
      Q => sig000000cb
    );
  blk000007d2 : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => sig00000773,
      R => sig000008b6,
      Q => NLW_blk000007d2_Q_UNCONNECTED
    );
  blk000007d3 : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => sig00000774,
      R => sig000008b6,
      Q => NLW_blk000007d3_Q_UNCONNECTED
    );
  blk000007d4 : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => sig00000775,
      R => sig000008b6,
      Q => NLW_blk000007d4_Q_UNCONNECTED
    );
  blk000007d5 : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => sig00000776,
      R => sig000008b6,
      Q => NLW_blk000007d5_Q_UNCONNECTED
    );
  blk000007d6 : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => sig00000777,
      R => sig000008b6,
      Q => NLW_blk000007d6_Q_UNCONNECTED
    );
  blk000007d7 : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => sig00000778,
      R => sig000008b6,
      Q => NLW_blk000007d7_Q_UNCONNECTED
    );
  blk000007d8 : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => sig00000779,
      R => sig000008b6,
      Q => NLW_blk000007d8_Q_UNCONNECTED
    );
  blk000007d9 : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => sig0000077a,
      R => sig000008b6,
      Q => NLW_blk000007d9_Q_UNCONNECTED
    );
  blk000007da : LUT6
    generic map(
      INIT => X"FF00F0F0CCCCAAAA"
    )
    port map (
      I0 => sig00000994,
      I1 => sig00000994,
      I2 => sig00000994,
      I3 => sig00000994,
      I4 => sig00000a59,
      I5 => sig00000a5a,
      O => sig00000764
    );
  blk000007db : LUT6
    generic map(
      INIT => X"FF00F0F0CCCCAAAA"
    )
    port map (
      I0 => sig00000993,
      I1 => sig00000994,
      I2 => sig00000994,
      I3 => sig00000994,
      I4 => sig00000a59,
      I5 => sig00000a5a,
      O => sig00000765
    );
  blk000007dc : LUT6
    generic map(
      INIT => X"FF00F0F0CCCCAAAA"
    )
    port map (
      I0 => sig00000992,
      I1 => sig00000993,
      I2 => sig00000994,
      I3 => sig00000994,
      I4 => sig00000a59,
      I5 => sig00000a5a,
      O => sig00000766
    );
  blk000007dd : LUT6
    generic map(
      INIT => X"FF00F0F0CCCCAAAA"
    )
    port map (
      I0 => sig00000991,
      I1 => sig00000992,
      I2 => sig00000993,
      I3 => sig00000994,
      I4 => sig00000a59,
      I5 => sig00000a5a,
      O => sig00000767
    );
  blk000007de : LUT6
    generic map(
      INIT => X"FF00F0F0CCCCAAAA"
    )
    port map (
      I0 => sig00000990,
      I1 => sig00000991,
      I2 => sig00000992,
      I3 => sig00000993,
      I4 => sig00000a59,
      I5 => sig00000a5a,
      O => sig00000768
    );
  blk000007df : LUT6
    generic map(
      INIT => X"FF00F0F0CCCCAAAA"
    )
    port map (
      I0 => sig0000098f,
      I1 => sig00000990,
      I2 => sig00000991,
      I3 => sig00000992,
      I4 => sig00000a59,
      I5 => sig00000a5a,
      O => sig00000769
    );
  blk000007e0 : LUT6
    generic map(
      INIT => X"FF00F0F0CCCCAAAA"
    )
    port map (
      I0 => sig0000098e,
      I1 => sig0000098f,
      I2 => sig00000990,
      I3 => sig00000991,
      I4 => sig00000a59,
      I5 => sig00000a5a,
      O => sig0000076a
    );
  blk000007e1 : LUT6
    generic map(
      INIT => X"FF00F0F0CCCCAAAA"
    )
    port map (
      I0 => sig0000098d,
      I1 => sig0000098e,
      I2 => sig0000098f,
      I3 => sig00000990,
      I4 => sig00000a59,
      I5 => sig00000a5a,
      O => sig0000076b
    );
  blk000007e2 : LUT6
    generic map(
      INIT => X"FF00F0F0CCCCAAAA"
    )
    port map (
      I0 => sig0000098c,
      I1 => sig0000098d,
      I2 => sig0000098e,
      I3 => sig0000098f,
      I4 => sig00000a59,
      I5 => sig00000a5a,
      O => sig0000076c
    );
  blk000007e3 : LUT6
    generic map(
      INIT => X"FF00F0F0CCCCAAAA"
    )
    port map (
      I0 => sig0000098b,
      I1 => sig0000098c,
      I2 => sig0000098d,
      I3 => sig0000098e,
      I4 => sig00000a59,
      I5 => sig00000a5a,
      O => sig0000076d
    );
  blk000007e4 : LUT6
    generic map(
      INIT => X"FF00F0F0CCCCAAAA"
    )
    port map (
      I0 => sig0000098a,
      I1 => sig0000098b,
      I2 => sig0000098c,
      I3 => sig0000098d,
      I4 => sig00000a59,
      I5 => sig00000a5a,
      O => sig0000076e
    );
  blk000007e5 : LUT6
    generic map(
      INIT => X"FF00F0F0CCCCAAAA"
    )
    port map (
      I0 => sig00000989,
      I1 => sig0000098a,
      I2 => sig0000098b,
      I3 => sig0000098c,
      I4 => sig00000a59,
      I5 => sig00000a5a,
      O => sig0000076f
    );
  blk000007e6 : LUT6
    generic map(
      INIT => X"FF00F0F0CCCCAAAA"
    )
    port map (
      I0 => sig00000988,
      I1 => sig00000989,
      I2 => sig0000098a,
      I3 => sig0000098b,
      I4 => sig00000a59,
      I5 => sig00000a5a,
      O => sig00000770
    );
  blk000007e7 : LUT6
    generic map(
      INIT => X"FF00F0F0CCCCAAAA"
    )
    port map (
      I0 => sig00000987,
      I1 => sig00000988,
      I2 => sig00000989,
      I3 => sig0000098a,
      I4 => sig00000a59,
      I5 => sig00000a5a,
      O => sig00000771
    );
  blk000007e8 : LUT6
    generic map(
      INIT => X"FF00F0F0CCCCAAAA"
    )
    port map (
      I0 => sig00000986,
      I1 => sig00000987,
      I2 => sig00000988,
      I3 => sig00000989,
      I4 => sig00000a59,
      I5 => sig00000a5a,
      O => sig00000772
    );
  blk000007e9 : LUT6
    generic map(
      INIT => X"FF00F0F0CCCCAAAA"
    )
    port map (
      I0 => sig00000985,
      I1 => sig00000986,
      I2 => sig00000987,
      I3 => sig00000988,
      I4 => sig00000a59,
      I5 => sig00000a5a,
      O => sig00000773
    );
  blk000007ea : LUT6
    generic map(
      INIT => X"FF00F0F0CCCCAAAA"
    )
    port map (
      I0 => sig00000984,
      I1 => sig00000985,
      I2 => sig00000986,
      I3 => sig00000987,
      I4 => sig00000a59,
      I5 => sig00000a5a,
      O => sig00000774
    );
  blk000007eb : LUT6
    generic map(
      INIT => X"FF00F0F0CCCCAAAA"
    )
    port map (
      I0 => sig00000983,
      I1 => sig00000984,
      I2 => sig00000985,
      I3 => sig00000986,
      I4 => sig00000a59,
      I5 => sig00000a5a,
      O => sig00000775
    );
  blk000007ec : LUT6
    generic map(
      INIT => X"FF00F0F0CCCCAAAA"
    )
    port map (
      I0 => sig00000982,
      I1 => sig00000983,
      I2 => sig00000984,
      I3 => sig00000985,
      I4 => sig00000a59,
      I5 => sig00000a5a,
      O => sig00000776
    );
  blk000007ed : LUT6
    generic map(
      INIT => X"FF00F0F0CCCCAAAA"
    )
    port map (
      I0 => sig00000981,
      I1 => sig00000982,
      I2 => sig00000983,
      I3 => sig00000984,
      I4 => sig00000a59,
      I5 => sig00000a5a,
      O => sig00000777
    );
  blk000007ee : LUT6
    generic map(
      INIT => X"FF00F0F0CCCCAAAA"
    )
    port map (
      I0 => sig000008b6,
      I1 => sig00000981,
      I2 => sig00000982,
      I3 => sig00000983,
      I4 => sig00000a59,
      I5 => sig00000a5a,
      O => sig00000778
    );
  blk000007ef : LUT6
    generic map(
      INIT => X"FF00F0F0CCCCAAAA"
    )
    port map (
      I0 => sig000008b6,
      I1 => sig000008b6,
      I2 => sig00000981,
      I3 => sig00000982,
      I4 => sig00000a59,
      I5 => sig00000a5a,
      O => sig00000779
    );
  blk000007f0 : LUT6
    generic map(
      INIT => X"FF00F0F0CCCCAAAA"
    )
    port map (
      I0 => sig000008b6,
      I1 => sig000008b6,
      I2 => sig000008b6,
      I3 => sig00000981,
      I4 => sig00000a59,
      I5 => sig00000a5a,
      O => sig0000077a
    );
  blk000007f1 : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => sig0000077b,
      R => sig000008b6,
      Q => NLW_blk000007f1_Q_UNCONNECTED
    );
  blk000007f2 : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => sig0000077c,
      R => sig000008b6,
      Q => NLW_blk000007f2_Q_UNCONNECTED
    );
  blk000007f3 : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => sig0000077d,
      R => sig000008b6,
      Q => NLW_blk000007f3_Q_UNCONNECTED
    );
  blk000007f4 : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => sig0000077e,
      R => sig000008b6,
      Q => sig000000e2
    );
  blk000007f5 : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => sig0000077f,
      R => sig000008b6,
      Q => sig000000e1
    );
  blk000007f6 : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => sig00000780,
      R => sig000008b6,
      Q => sig000000e0
    );
  blk000007f7 : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => sig00000781,
      R => sig000008b6,
      Q => sig000000df
    );
  blk000007f8 : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => sig00000782,
      R => sig000008b6,
      Q => sig000000de
    );
  blk000007f9 : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => sig00000783,
      R => sig000008b6,
      Q => sig000000dd
    );
  blk000007fa : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => sig00000784,
      R => sig000008b6,
      Q => sig000000dc
    );
  blk000007fb : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => sig00000785,
      R => sig000008b6,
      Q => sig000000db
    );
  blk000007fc : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => sig00000786,
      R => sig000008b6,
      Q => sig000000da
    );
  blk000007fd : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => sig00000787,
      R => sig000008b6,
      Q => sig000000d9
    );
  blk000007fe : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => sig00000788,
      R => sig000008b6,
      Q => sig000000d8
    );
  blk000007ff : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => sig00000789,
      R => sig000008b6,
      Q => sig000000d7
    );
  blk00000800 : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => sig0000078a,
      R => sig000008b6,
      Q => NLW_blk00000800_Q_UNCONNECTED
    );
  blk00000801 : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => sig0000078b,
      R => sig000008b6,
      Q => NLW_blk00000801_Q_UNCONNECTED
    );
  blk00000802 : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => sig0000078c,
      R => sig000008b6,
      Q => NLW_blk00000802_Q_UNCONNECTED
    );
  blk00000803 : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => sig0000078d,
      R => sig000008b6,
      Q => NLW_blk00000803_Q_UNCONNECTED
    );
  blk00000804 : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => sig0000078e,
      R => sig000008b6,
      Q => NLW_blk00000804_Q_UNCONNECTED
    );
  blk00000805 : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => sig0000078f,
      R => sig000008b6,
      Q => NLW_blk00000805_Q_UNCONNECTED
    );
  blk00000806 : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => sig00000790,
      R => sig000008b6,
      Q => NLW_blk00000806_Q_UNCONNECTED
    );
  blk00000807 : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => sig00000791,
      R => sig000008b6,
      Q => NLW_blk00000807_Q_UNCONNECTED
    );
  blk00000808 : LUT6
    generic map(
      INIT => X"FF00F0F0CCCCAAAA"
    )
    port map (
      I0 => sig000008e8,
      I1 => sig000008e8,
      I2 => sig000008e8,
      I3 => sig000008e8,
      I4 => sig00000a59,
      I5 => sig00000a5a,
      O => sig0000077b
    );
  blk00000809 : LUT6
    generic map(
      INIT => X"FF00F0F0CCCCAAAA"
    )
    port map (
      I0 => sig000008e7,
      I1 => sig000008e8,
      I2 => sig000008e8,
      I3 => sig000008e8,
      I4 => sig00000a59,
      I5 => sig00000a5a,
      O => sig0000077c
    );
  blk0000080a : LUT6
    generic map(
      INIT => X"FF00F0F0CCCCAAAA"
    )
    port map (
      I0 => sig000008e6,
      I1 => sig000008e7,
      I2 => sig000008e8,
      I3 => sig000008e8,
      I4 => sig00000a59,
      I5 => sig00000a5a,
      O => sig0000077d
    );
  blk0000080b : LUT6
    generic map(
      INIT => X"FF00F0F0CCCCAAAA"
    )
    port map (
      I0 => sig000008e5,
      I1 => sig000008e6,
      I2 => sig000008e7,
      I3 => sig000008e8,
      I4 => sig00000a59,
      I5 => sig00000a5a,
      O => sig0000077e
    );
  blk0000080c : LUT6
    generic map(
      INIT => X"FF00F0F0CCCCAAAA"
    )
    port map (
      I0 => sig000008e4,
      I1 => sig000008e5,
      I2 => sig000008e6,
      I3 => sig000008e7,
      I4 => sig00000a59,
      I5 => sig00000a5a,
      O => sig0000077f
    );
  blk0000080d : LUT6
    generic map(
      INIT => X"FF00F0F0CCCCAAAA"
    )
    port map (
      I0 => sig000008e3,
      I1 => sig000008e4,
      I2 => sig000008e5,
      I3 => sig000008e6,
      I4 => sig00000a59,
      I5 => sig00000a5a,
      O => sig00000780
    );
  blk0000080e : LUT6
    generic map(
      INIT => X"FF00F0F0CCCCAAAA"
    )
    port map (
      I0 => sig000008e2,
      I1 => sig000008e3,
      I2 => sig000008e4,
      I3 => sig000008e5,
      I4 => sig00000a59,
      I5 => sig00000a5a,
      O => sig00000781
    );
  blk0000080f : LUT6
    generic map(
      INIT => X"FF00F0F0CCCCAAAA"
    )
    port map (
      I0 => sig000008e1,
      I1 => sig000008e2,
      I2 => sig000008e3,
      I3 => sig000008e4,
      I4 => sig00000a59,
      I5 => sig00000a5a,
      O => sig00000782
    );
  blk00000810 : LUT6
    generic map(
      INIT => X"FF00F0F0CCCCAAAA"
    )
    port map (
      I0 => sig000008e0,
      I1 => sig000008e1,
      I2 => sig000008e2,
      I3 => sig000008e3,
      I4 => sig00000a59,
      I5 => sig00000a5a,
      O => sig00000783
    );
  blk00000811 : LUT6
    generic map(
      INIT => X"FF00F0F0CCCCAAAA"
    )
    port map (
      I0 => sig000008df,
      I1 => sig000008e0,
      I2 => sig000008e1,
      I3 => sig000008e2,
      I4 => sig00000a59,
      I5 => sig00000a5a,
      O => sig00000784
    );
  blk00000812 : LUT6
    generic map(
      INIT => X"FF00F0F0CCCCAAAA"
    )
    port map (
      I0 => sig000008de,
      I1 => sig000008df,
      I2 => sig000008e0,
      I3 => sig000008e1,
      I4 => sig00000a59,
      I5 => sig00000a5a,
      O => sig00000785
    );
  blk00000813 : LUT6
    generic map(
      INIT => X"FF00F0F0CCCCAAAA"
    )
    port map (
      I0 => sig000008dd,
      I1 => sig000008de,
      I2 => sig000008df,
      I3 => sig000008e0,
      I4 => sig00000a59,
      I5 => sig00000a5a,
      O => sig00000786
    );
  blk00000814 : LUT6
    generic map(
      INIT => X"FF00F0F0CCCCAAAA"
    )
    port map (
      I0 => sig000008dc,
      I1 => sig000008dd,
      I2 => sig000008de,
      I3 => sig000008df,
      I4 => sig00000a59,
      I5 => sig00000a5a,
      O => sig00000787
    );
  blk00000815 : LUT6
    generic map(
      INIT => X"FF00F0F0CCCCAAAA"
    )
    port map (
      I0 => sig000008db,
      I1 => sig000008dc,
      I2 => sig000008dd,
      I3 => sig000008de,
      I4 => sig00000a59,
      I5 => sig00000a5a,
      O => sig00000788
    );
  blk00000816 : LUT6
    generic map(
      INIT => X"FF00F0F0CCCCAAAA"
    )
    port map (
      I0 => sig000008da,
      I1 => sig000008db,
      I2 => sig000008dc,
      I3 => sig000008dd,
      I4 => sig00000a59,
      I5 => sig00000a5a,
      O => sig00000789
    );
  blk00000817 : LUT6
    generic map(
      INIT => X"FF00F0F0CCCCAAAA"
    )
    port map (
      I0 => sig000008d9,
      I1 => sig000008da,
      I2 => sig000008db,
      I3 => sig000008dc,
      I4 => sig00000a59,
      I5 => sig00000a5a,
      O => sig0000078a
    );
  blk00000818 : LUT6
    generic map(
      INIT => X"FF00F0F0CCCCAAAA"
    )
    port map (
      I0 => sig000008d8,
      I1 => sig000008d9,
      I2 => sig000008da,
      I3 => sig000008db,
      I4 => sig00000a59,
      I5 => sig00000a5a,
      O => sig0000078b
    );
  blk00000819 : LUT6
    generic map(
      INIT => X"FF00F0F0CCCCAAAA"
    )
    port map (
      I0 => sig000008d7,
      I1 => sig000008d8,
      I2 => sig000008d9,
      I3 => sig000008da,
      I4 => sig00000a59,
      I5 => sig00000a5a,
      O => sig0000078c
    );
  blk0000081a : LUT6
    generic map(
      INIT => X"FF00F0F0CCCCAAAA"
    )
    port map (
      I0 => sig000008d6,
      I1 => sig000008d7,
      I2 => sig000008d8,
      I3 => sig000008d9,
      I4 => sig00000a59,
      I5 => sig00000a5a,
      O => sig0000078d
    );
  blk0000081b : LUT6
    generic map(
      INIT => X"FF00F0F0CCCCAAAA"
    )
    port map (
      I0 => sig000008d5,
      I1 => sig000008d6,
      I2 => sig000008d7,
      I3 => sig000008d8,
      I4 => sig00000a59,
      I5 => sig00000a5a,
      O => sig0000078e
    );
  blk0000081c : LUT6
    generic map(
      INIT => X"FF00F0F0CCCCAAAA"
    )
    port map (
      I0 => sig000008b6,
      I1 => sig000008d5,
      I2 => sig000008d6,
      I3 => sig000008d7,
      I4 => sig00000a59,
      I5 => sig00000a5a,
      O => sig0000078f
    );
  blk0000081d : LUT6
    generic map(
      INIT => X"FF00F0F0CCCCAAAA"
    )
    port map (
      I0 => sig000008b6,
      I1 => sig000008b6,
      I2 => sig000008d5,
      I3 => sig000008d6,
      I4 => sig00000a59,
      I5 => sig00000a5a,
      O => sig00000790
    );
  blk0000081e : LUT6
    generic map(
      INIT => X"FF00F0F0CCCCAAAA"
    )
    port map (
      I0 => sig000008b6,
      I1 => sig000008b6,
      I2 => sig000008b6,
      I3 => sig000008d5,
      I4 => sig00000a59,
      I5 => sig00000a5a,
      O => sig00000791
    );
  blk00000828 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => sig0000087a,
      Q => sig0000080d
    );
  blk00000829 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => sig00000879,
      Q => sig0000080c
    );
  blk0000082a : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => sig00000878,
      Q => sig0000080b
    );
  blk0000082b : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => sig00000877,
      Q => sig0000080a
    );
  blk0000082c : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => sig00000876,
      Q => sig00000851
    );
  blk0000082d : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => sig00000875,
      Q => sig00000850
    );
  blk0000082e : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => sig00000874,
      Q => sig0000084f
    );
  blk0000082f : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => sig00000873,
      Q => sig0000084e
    );
  blk00000830 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => sig00000a49,
      Q => sig00000831
    );
  blk00000831 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => sig00000a4a,
      Q => sig00000830
    );
  blk00000832 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => sig00000a4b,
      Q => sig0000082f
    );
  blk00000833 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => sig00000a4c,
      Q => sig0000082e
    );
  blk00000834 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => sig00000a4d,
      Q => sig0000082d
    );
  blk00000835 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => sig00000a4e,
      Q => sig0000082c
    );
  blk00000836 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => sig00000a4f,
      Q => sig0000082b
    );
  blk00000837 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => sig00000a50,
      Q => sig0000082a
    );
  blk00000838 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => sig00000a51,
      Q => sig00000829
    );
  blk00000839 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => sig00000a52,
      Q => sig00000828
    );
  blk0000083a : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => sig00000a53,
      Q => sig00000827
    );
  blk0000083b : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => sig00000a54,
      Q => sig00000826
    );
  blk0000083c : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => sig00000a55,
      Q => sig00000825
    );
  blk0000083d : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => sig00000a56,
      Q => sig00000824
    );
  blk0000083e : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => sig00000a3b,
      Q => sig000007f3
    );
  blk0000083f : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => sig00000a3c,
      Q => sig000007f2
    );
  blk00000840 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => sig00000a3d,
      Q => sig000007f1
    );
  blk00000841 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => sig00000a3e,
      Q => sig000007f0
    );
  blk00000842 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => sig00000a3f,
      Q => sig000007ef
    );
  blk00000843 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => sig00000a40,
      Q => sig000007ee
    );
  blk00000844 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => sig00000a41,
      Q => sig000007ed
    );
  blk00000845 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => sig00000a42,
      Q => sig000007ec
    );
  blk00000846 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => sig00000a43,
      Q => sig000007eb
    );
  blk00000847 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => sig00000a44,
      Q => sig000007ea
    );
  blk00000848 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => sig00000a45,
      Q => sig000007e9
    );
  blk00000849 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => sig00000a46,
      Q => sig000007e8
    );
  blk0000084a : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => sig00000a47,
      Q => sig000007e7
    );
  blk0000084b : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => sig00000a48,
      Q => sig000007e6
    );
  blk0000084c : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => sig000007bd,
      Q => sig00000809
    );
  blk0000084d : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => sig000007bc,
      Q => sig00000808
    );
  blk0000084e : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => sig000007bb,
      Q => sig00000807
    );
  blk0000084f : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => sig000007ba,
      Q => sig00000806
    );
  blk00000850 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => sig000007b9,
      Q => sig00000805
    );
  blk00000851 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => sig000007b8,
      Q => sig00000804
    );
  blk00000852 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => sig000007b7,
      Q => sig00000803
    );
  blk00000853 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => sig000007b6,
      Q => sig00000802
    );
  blk00000854 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => sig000007b5,
      Q => sig00000801
    );
  blk00000855 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => sig000007b4,
      Q => sig00000800
    );
  blk00000856 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => sig000007b3,
      Q => sig000007ff
    );
  blk00000857 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => sig000007a7,
      Q => sig000007fe
    );
  blk00000858 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => sig000007a6,
      Q => sig000007fd
    );
  blk00000859 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => sig000007a5,
      Q => sig000007fc
    );
  blk0000085a : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => sig000007a4,
      Q => sig000007fb
    );
  blk0000085b : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => sig000007a3,
      Q => sig000007fa
    );
  blk0000085c : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => sig000007a2,
      Q => sig000007f9
    );
  blk0000085d : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => sig000007a1,
      Q => sig000007f8
    );
  blk0000085e : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => sig000007a0,
      Q => sig000007f7
    );
  blk0000085f : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => sig0000079f,
      Q => sig000007f6
    );
  blk00000860 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => sig0000079e,
      Q => sig000007f5
    );
  blk00000861 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => sig0000079d,
      Q => sig000007f4
    );
  blk00000862 : MUXCY
    port map (
      CI => sig000006d1,
      DI => sig000008b6,
      S => sig000007be,
      O => sig000007bf
    );
  blk00000863 : XORCY
    port map (
      CI => sig000006d1,
      LI => sig000007be,
      O => sig0000079c
    );
  blk00000864 : MUXCY
    port map (
      CI => sig000007bf,
      DI => sig000008b6,
      S => sig000007c0,
      O => sig000007c1
    );
  blk00000865 : XORCY
    port map (
      CI => sig000007bf,
      LI => sig000007c0,
      O => sig0000079b
    );
  blk00000866 : MUXCY
    port map (
      CI => sig000007c1,
      DI => sig000008b6,
      S => sig000007c2,
      O => sig000007c3
    );
  blk00000867 : XORCY
    port map (
      CI => sig000007c1,
      LI => sig000007c2,
      O => sig0000079a
    );
  blk00000868 : MUXCY
    port map (
      CI => sig000007c3,
      DI => sig000008b6,
      S => sig000007c4,
      O => sig000007c5
    );
  blk00000869 : XORCY
    port map (
      CI => sig000007c3,
      LI => sig000007c4,
      O => sig00000799
    );
  blk0000086a : MUXCY
    port map (
      CI => sig000007c5,
      DI => sig000008b6,
      S => sig000007c6,
      O => sig000007c7
    );
  blk0000086b : XORCY
    port map (
      CI => sig000007c5,
      LI => sig000007c6,
      O => sig00000798
    );
  blk0000086c : MUXCY
    port map (
      CI => sig000007c7,
      DI => sig000008b6,
      S => sig000007c8,
      O => sig000007c9
    );
  blk0000086d : XORCY
    port map (
      CI => sig000007c7,
      LI => sig000007c8,
      O => sig00000797
    );
  blk0000086e : MUXCY
    port map (
      CI => sig000007c9,
      DI => sig000008b6,
      S => sig000007ca,
      O => sig000007cb
    );
  blk0000086f : XORCY
    port map (
      CI => sig000007c9,
      LI => sig000007ca,
      O => sig00000796
    );
  blk00000870 : MUXCY
    port map (
      CI => sig000007cb,
      DI => sig000008b6,
      S => sig000007cc,
      O => sig000007cd
    );
  blk00000871 : XORCY
    port map (
      CI => sig000007cb,
      LI => sig000007cc,
      O => sig00000795
    );
  blk00000872 : MUXCY
    port map (
      CI => sig000007cd,
      DI => sig000008b6,
      S => sig000007ce,
      O => sig000007cf
    );
  blk00000873 : XORCY
    port map (
      CI => sig000007cd,
      LI => sig000007ce,
      O => sig00000794
    );
  blk00000874 : MUXCY
    port map (
      CI => sig000007cf,
      DI => sig000008b6,
      S => sig000007d0,
      O => sig000007d1
    );
  blk00000875 : XORCY
    port map (
      CI => sig000007cf,
      LI => sig000007d0,
      O => sig00000793
    );
  blk00000876 : XORCY
    port map (
      CI => sig000007d1,
      LI => sig000006d1,
      O => sig00000792
    );
  blk00000877 : MUXCY
    port map (
      CI => sig000006d1,
      DI => sig000008b6,
      S => sig000007d2,
      O => sig000007d3
    );
  blk00000878 : XORCY
    port map (
      CI => sig000006d1,
      LI => sig000007d2,
      O => sig000007b2
    );
  blk00000879 : MUXCY
    port map (
      CI => sig000007d3,
      DI => sig000008b6,
      S => sig000007d4,
      O => sig000007d5
    );
  blk0000087a : XORCY
    port map (
      CI => sig000007d3,
      LI => sig000007d4,
      O => sig000007b1
    );
  blk0000087b : MUXCY
    port map (
      CI => sig000007d5,
      DI => sig000008b6,
      S => sig000007d6,
      O => sig000007d7
    );
  blk0000087c : XORCY
    port map (
      CI => sig000007d5,
      LI => sig000007d6,
      O => sig000007b0
    );
  blk0000087d : MUXCY
    port map (
      CI => sig000007d7,
      DI => sig000008b6,
      S => sig000007d8,
      O => sig000007d9
    );
  blk0000087e : XORCY
    port map (
      CI => sig000007d7,
      LI => sig000007d8,
      O => sig000007af
    );
  blk0000087f : MUXCY
    port map (
      CI => sig000007d9,
      DI => sig000008b6,
      S => sig000007da,
      O => sig000007db
    );
  blk00000880 : XORCY
    port map (
      CI => sig000007d9,
      LI => sig000007da,
      O => sig000007ae
    );
  blk00000881 : MUXCY
    port map (
      CI => sig000007db,
      DI => sig000008b6,
      S => sig000007dc,
      O => sig000007dd
    );
  blk00000882 : XORCY
    port map (
      CI => sig000007db,
      LI => sig000007dc,
      O => sig000007ad
    );
  blk00000883 : MUXCY
    port map (
      CI => sig000007dd,
      DI => sig000008b6,
      S => sig000007de,
      O => sig000007df
    );
  blk00000884 : XORCY
    port map (
      CI => sig000007dd,
      LI => sig000007de,
      O => sig000007ac
    );
  blk00000885 : MUXCY
    port map (
      CI => sig000007df,
      DI => sig000008b6,
      S => sig000007e0,
      O => sig000007e1
    );
  blk00000886 : XORCY
    port map (
      CI => sig000007df,
      LI => sig000007e0,
      O => sig000007ab
    );
  blk00000887 : MUXCY
    port map (
      CI => sig000007e1,
      DI => sig000008b6,
      S => sig000007e2,
      O => sig000007e3
    );
  blk00000888 : XORCY
    port map (
      CI => sig000007e1,
      LI => sig000007e2,
      O => sig000007aa
    );
  blk00000889 : MUXCY
    port map (
      CI => sig000007e3,
      DI => sig000008b6,
      S => sig000007e4,
      O => sig000007e5
    );
  blk0000088a : XORCY
    port map (
      CI => sig000007e3,
      LI => sig000007e4,
      O => sig000007a9
    );
  blk0000088b : XORCY
    port map (
      CI => sig000007e5,
      LI => sig000006d1,
      O => sig000007a8
    );
  blk0000088c : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => sig000008a3,
      Q => sig00000872
    );
  blk0000088d : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => sig000008a2,
      Q => sig00000871
    );
  blk0000088e : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => sig000008a1,
      Q => sig00000870
    );
  blk0000088f : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => sig000008a0,
      Q => sig0000086f
    );
  blk00000890 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => sig0000089f,
      Q => sig0000086e
    );
  blk00000891 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => sig0000089e,
      Q => sig0000086d
    );
  blk00000892 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => sig0000089d,
      Q => sig0000086c
    );
  blk00000893 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => sig0000089c,
      Q => sig0000086b
    );
  blk00000894 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => sig0000089b,
      Q => sig0000086a
    );
  blk00000895 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => sig0000089a,
      Q => sig00000869
    );
  blk00000896 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => sig00000899,
      Q => sig00000868
    );
  blk00000897 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => sig00000898,
      Q => sig00000867
    );
  blk00000898 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => sig0000088c,
      Q => sig00000876
    );
  blk00000899 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => sig0000088b,
      Q => sig00000875
    );
  blk0000089a : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => sig0000088a,
      Q => sig00000874
    );
  blk0000089b : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => sig00000889,
      Q => sig00000873
    );
  blk0000089c : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => sig0000087e,
      Q => sig0000087a
    );
  blk0000089d : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => sig0000087d,
      Q => sig00000879
    );
  blk0000089e : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => sig0000087c,
      Q => sig00000878
    );
  blk0000089f : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => sig0000087b,
      Q => sig00000877
    );
  blk000008a0 : LUT2
    generic map(
      INIT => X"6"
    )
    port map (
      I0 => sig000007fe,
      I1 => sig00000809,
      O => sig000009a7
    );
  blk000008a1 : MUXCY
    port map (
      CI => sig000008b6,
      DI => sig000007fe,
      S => sig000009a7,
      O => sig000009a8
    );
  blk000008a2 : XORCY
    port map (
      CI => sig000008b6,
      LI => sig000009a7,
      O => sig000008a3
    );
  blk000008a3 : LUT2
    generic map(
      INIT => X"6"
    )
    port map (
      I0 => sig000007fd,
      I1 => sig00000808,
      O => sig000009a9
    );
  blk000008a4 : MUXCY
    port map (
      CI => sig000009a8,
      DI => sig000007fd,
      S => sig000009a9,
      O => sig000009aa
    );
  blk000008a5 : XORCY
    port map (
      CI => sig000009a8,
      LI => sig000009a9,
      O => sig000008a2
    );
  blk000008a6 : LUT2
    generic map(
      INIT => X"6"
    )
    port map (
      I0 => sig000007fc,
      I1 => sig00000807,
      O => sig000009ab
    );
  blk000008a7 : MUXCY
    port map (
      CI => sig000009aa,
      DI => sig000007fc,
      S => sig000009ab,
      O => sig000009ac
    );
  blk000008a8 : XORCY
    port map (
      CI => sig000009aa,
      LI => sig000009ab,
      O => sig000008a1
    );
  blk000008a9 : LUT2
    generic map(
      INIT => X"6"
    )
    port map (
      I0 => sig000007fb,
      I1 => sig00000806,
      O => sig000009ad
    );
  blk000008aa : MUXCY
    port map (
      CI => sig000009ac,
      DI => sig000007fb,
      S => sig000009ad,
      O => sig000009ae
    );
  blk000008ab : XORCY
    port map (
      CI => sig000009ac,
      LI => sig000009ad,
      O => sig000008a0
    );
  blk000008ac : LUT2
    generic map(
      INIT => X"6"
    )
    port map (
      I0 => sig000007fa,
      I1 => sig00000805,
      O => sig000009af
    );
  blk000008ad : MUXCY
    port map (
      CI => sig000009ae,
      DI => sig000007fa,
      S => sig000009af,
      O => sig000009b0
    );
  blk000008ae : XORCY
    port map (
      CI => sig000009ae,
      LI => sig000009af,
      O => sig0000089f
    );
  blk000008af : LUT2
    generic map(
      INIT => X"6"
    )
    port map (
      I0 => sig000007f9,
      I1 => sig00000804,
      O => sig000009b1
    );
  blk000008b0 : MUXCY
    port map (
      CI => sig000009b0,
      DI => sig000007f9,
      S => sig000009b1,
      O => sig000009b2
    );
  blk000008b1 : XORCY
    port map (
      CI => sig000009b0,
      LI => sig000009b1,
      O => sig0000089e
    );
  blk000008b2 : LUT2
    generic map(
      INIT => X"6"
    )
    port map (
      I0 => sig000007f8,
      I1 => sig00000803,
      O => sig000009b3
    );
  blk000008b3 : MUXCY
    port map (
      CI => sig000009b2,
      DI => sig000007f8,
      S => sig000009b3,
      O => sig000009b4
    );
  blk000008b4 : XORCY
    port map (
      CI => sig000009b2,
      LI => sig000009b3,
      O => sig0000089d
    );
  blk000008b5 : LUT2
    generic map(
      INIT => X"6"
    )
    port map (
      I0 => sig000007f7,
      I1 => sig00000802,
      O => sig000009b5
    );
  blk000008b6 : MUXCY
    port map (
      CI => sig000009b4,
      DI => sig000007f7,
      S => sig000009b5,
      O => sig000009b6
    );
  blk000008b7 : XORCY
    port map (
      CI => sig000009b4,
      LI => sig000009b5,
      O => sig0000089c
    );
  blk000008b8 : LUT2
    generic map(
      INIT => X"6"
    )
    port map (
      I0 => sig000007f6,
      I1 => sig00000801,
      O => sig000009b7
    );
  blk000008b9 : MUXCY
    port map (
      CI => sig000009b6,
      DI => sig000007f6,
      S => sig000009b7,
      O => sig000009b8
    );
  blk000008ba : XORCY
    port map (
      CI => sig000009b6,
      LI => sig000009b7,
      O => sig0000089b
    );
  blk000008bb : LUT2
    generic map(
      INIT => X"6"
    )
    port map (
      I0 => sig000007f5,
      I1 => sig00000800,
      O => sig000009b9
    );
  blk000008bc : MUXCY
    port map (
      CI => sig000009b8,
      DI => sig000007f5,
      S => sig000009b9,
      O => sig000009ba
    );
  blk000008bd : XORCY
    port map (
      CI => sig000009b8,
      LI => sig000009b9,
      O => sig0000089a
    );
  blk000008be : LUT2
    generic map(
      INIT => X"6"
    )
    port map (
      I0 => sig000007f4,
      I1 => sig000007ff,
      O => sig000009bb
    );
  blk000008bf : MUXCY
    port map (
      CI => sig000009ba,
      DI => sig000007f4,
      S => sig00000ef0,
      O => sig000009bc
    );
  blk000008c0 : XORCY
    port map (
      CI => sig000009ba,
      LI => sig00000ef0,
      O => sig00000899
    );
  blk000008c1 : XORCY
    port map (
      CI => sig000009bc,
      LI => sig000009bb,
      O => sig00000898
    );
  blk000008c2 : LUT2
    generic map(
      INIT => X"6"
    )
    port map (
      I0 => sig00000831,
      I1 => sig000007f3,
      O => sig000009bd
    );
  blk000008c3 : MUXCY
    port map (
      CI => sig000008b6,
      DI => sig00000831,
      S => sig000009bd,
      O => sig000009be
    );
  blk000008c4 : LUT2
    generic map(
      INIT => X"6"
    )
    port map (
      I0 => sig00000830,
      I1 => sig000007f2,
      O => sig000009bf
    );
  blk000008c5 : MUXCY
    port map (
      CI => sig000009be,
      DI => sig00000830,
      S => sig000009bf,
      O => sig000009c0
    );
  blk000008c6 : XORCY
    port map (
      CI => sig000009be,
      LI => sig000009bf,
      O => sig00000888
    );
  blk000008c7 : LUT2
    generic map(
      INIT => X"6"
    )
    port map (
      I0 => sig0000082f,
      I1 => sig000007f1,
      O => sig000009c1
    );
  blk000008c8 : MUXCY
    port map (
      CI => sig000009c0,
      DI => sig0000082f,
      S => sig000009c1,
      O => sig000009c2
    );
  blk000008c9 : XORCY
    port map (
      CI => sig000009c0,
      LI => sig000009c1,
      O => sig00000887
    );
  blk000008ca : LUT2
    generic map(
      INIT => X"6"
    )
    port map (
      I0 => sig0000082e,
      I1 => sig000007f0,
      O => sig000009c3
    );
  blk000008cb : MUXCY
    port map (
      CI => sig000009c2,
      DI => sig0000082e,
      S => sig000009c3,
      O => sig000009c4
    );
  blk000008cc : XORCY
    port map (
      CI => sig000009c2,
      LI => sig000009c3,
      O => sig00000886
    );
  blk000008cd : LUT2
    generic map(
      INIT => X"6"
    )
    port map (
      I0 => sig0000082d,
      I1 => sig000007ef,
      O => sig000009c5
    );
  blk000008ce : MUXCY
    port map (
      CI => sig000009c4,
      DI => sig0000082d,
      S => sig000009c5,
      O => sig000009c6
    );
  blk000008cf : XORCY
    port map (
      CI => sig000009c4,
      LI => sig000009c5,
      O => sig00000885
    );
  blk000008d0 : LUT2
    generic map(
      INIT => X"6"
    )
    port map (
      I0 => sig0000082c,
      I1 => sig000007ee,
      O => sig000009c7
    );
  blk000008d1 : MUXCY
    port map (
      CI => sig000009c6,
      DI => sig0000082c,
      S => sig000009c7,
      O => sig000009c8
    );
  blk000008d2 : XORCY
    port map (
      CI => sig000009c6,
      LI => sig000009c7,
      O => sig00000884
    );
  blk000008d3 : LUT2
    generic map(
      INIT => X"6"
    )
    port map (
      I0 => sig0000082b,
      I1 => sig000007ed,
      O => sig000009c9
    );
  blk000008d4 : MUXCY
    port map (
      CI => sig000009c8,
      DI => sig0000082b,
      S => sig000009c9,
      O => sig000009ca
    );
  blk000008d5 : XORCY
    port map (
      CI => sig000009c8,
      LI => sig000009c9,
      O => sig00000883
    );
  blk000008d6 : LUT2
    generic map(
      INIT => X"6"
    )
    port map (
      I0 => sig0000082a,
      I1 => sig000007ec,
      O => sig000009cb
    );
  blk000008d7 : MUXCY
    port map (
      CI => sig000009ca,
      DI => sig0000082a,
      S => sig000009cb,
      O => sig000009cc
    );
  blk000008d8 : XORCY
    port map (
      CI => sig000009ca,
      LI => sig000009cb,
      O => sig00000882
    );
  blk000008d9 : LUT2
    generic map(
      INIT => X"6"
    )
    port map (
      I0 => sig00000829,
      I1 => sig000007eb,
      O => sig000009cd
    );
  blk000008da : MUXCY
    port map (
      CI => sig000009cc,
      DI => sig00000829,
      S => sig000009cd,
      O => sig000009ce
    );
  blk000008db : XORCY
    port map (
      CI => sig000009cc,
      LI => sig000009cd,
      O => sig00000881
    );
  blk000008dc : LUT2
    generic map(
      INIT => X"6"
    )
    port map (
      I0 => sig00000828,
      I1 => sig000007ea,
      O => sig000009cf
    );
  blk000008dd : MUXCY
    port map (
      CI => sig000009ce,
      DI => sig00000828,
      S => sig000009cf,
      O => sig000009d0
    );
  blk000008de : XORCY
    port map (
      CI => sig000009ce,
      LI => sig000009cf,
      O => sig00000880
    );
  blk000008df : LUT2
    generic map(
      INIT => X"6"
    )
    port map (
      I0 => sig00000827,
      I1 => sig000007e9,
      O => sig000009d1
    );
  blk000008e0 : MUXCY
    port map (
      CI => sig000009d0,
      DI => sig00000827,
      S => sig000009d1,
      O => sig000009d2
    );
  blk000008e1 : XORCY
    port map (
      CI => sig000009d0,
      LI => sig000009d1,
      O => sig0000087f
    );
  blk000008e2 : LUT2
    generic map(
      INIT => X"6"
    )
    port map (
      I0 => sig00000826,
      I1 => sig000007e8,
      O => sig000009d3
    );
  blk000008e3 : MUXCY
    port map (
      CI => sig000009d2,
      DI => sig00000826,
      S => sig000009d3,
      O => sig000009d4
    );
  blk000008e4 : XORCY
    port map (
      CI => sig000009d2,
      LI => sig000009d3,
      O => sig0000087e
    );
  blk000008e5 : LUT2
    generic map(
      INIT => X"6"
    )
    port map (
      I0 => sig00000825,
      I1 => sig000007e7,
      O => sig000009d5
    );
  blk000008e6 : MUXCY
    port map (
      CI => sig000009d4,
      DI => sig00000825,
      S => sig000009d5,
      O => sig000009d6
    );
  blk000008e7 : XORCY
    port map (
      CI => sig000009d4,
      LI => sig000009d5,
      O => sig0000087d
    );
  blk000008e8 : LUT2
    generic map(
      INIT => X"6"
    )
    port map (
      I0 => sig00000824,
      I1 => sig000007e6,
      O => sig000009d7
    );
  blk000008e9 : MUXCY
    port map (
      CI => sig000009d6,
      DI => sig00000824,
      S => sig00000ef1,
      O => sig000009d8
    );
  blk000008ea : XORCY
    port map (
      CI => sig000009d6,
      LI => sig00000ef1,
      O => sig0000087c
    );
  blk000008eb : XORCY
    port map (
      CI => sig000009d8,
      LI => sig000009d7,
      O => sig0000087b
    );
  blk000008ec : LUT2
    generic map(
      INIT => X"9"
    )
    port map (
      I0 => sig000007f3,
      I1 => sig00000831,
      O => sig000009d9
    );
  blk000008ed : MUXCY
    port map (
      CI => sig000006d1,
      DI => sig000007f3,
      S => sig000009d9,
      O => sig000009da
    );
  blk000008ee : XORCY
    port map (
      CI => sig000006d1,
      LI => sig000009d9,
      O => sig00000897
    );
  blk000008ef : LUT2
    generic map(
      INIT => X"9"
    )
    port map (
      I0 => sig000007f2,
      I1 => sig00000830,
      O => sig000009db
    );
  blk000008f0 : MUXCY
    port map (
      CI => sig000009da,
      DI => sig000007f2,
      S => sig000009db,
      O => sig000009dc
    );
  blk000008f1 : XORCY
    port map (
      CI => sig000009da,
      LI => sig000009db,
      O => sig00000896
    );
  blk000008f2 : LUT2
    generic map(
      INIT => X"9"
    )
    port map (
      I0 => sig000007f1,
      I1 => sig0000082f,
      O => sig000009dd
    );
  blk000008f3 : MUXCY
    port map (
      CI => sig000009dc,
      DI => sig000007f1,
      S => sig000009dd,
      O => sig000009de
    );
  blk000008f4 : XORCY
    port map (
      CI => sig000009dc,
      LI => sig000009dd,
      O => sig00000895
    );
  blk000008f5 : LUT2
    generic map(
      INIT => X"9"
    )
    port map (
      I0 => sig000007f0,
      I1 => sig0000082e,
      O => sig000009df
    );
  blk000008f6 : MUXCY
    port map (
      CI => sig000009de,
      DI => sig000007f0,
      S => sig000009df,
      O => sig000009e0
    );
  blk000008f7 : XORCY
    port map (
      CI => sig000009de,
      LI => sig000009df,
      O => sig00000894
    );
  blk000008f8 : LUT2
    generic map(
      INIT => X"9"
    )
    port map (
      I0 => sig000007ef,
      I1 => sig0000082d,
      O => sig000009e1
    );
  blk000008f9 : MUXCY
    port map (
      CI => sig000009e0,
      DI => sig000007ef,
      S => sig000009e1,
      O => sig000009e2
    );
  blk000008fa : XORCY
    port map (
      CI => sig000009e0,
      LI => sig000009e1,
      O => sig00000893
    );
  blk000008fb : LUT2
    generic map(
      INIT => X"9"
    )
    port map (
      I0 => sig000007ee,
      I1 => sig0000082c,
      O => sig000009e3
    );
  blk000008fc : MUXCY
    port map (
      CI => sig000009e2,
      DI => sig000007ee,
      S => sig000009e3,
      O => sig000009e4
    );
  blk000008fd : XORCY
    port map (
      CI => sig000009e2,
      LI => sig000009e3,
      O => sig00000892
    );
  blk000008fe : LUT2
    generic map(
      INIT => X"9"
    )
    port map (
      I0 => sig000007ed,
      I1 => sig0000082b,
      O => sig000009e5
    );
  blk000008ff : MUXCY
    port map (
      CI => sig000009e4,
      DI => sig000007ed,
      S => sig000009e5,
      O => sig000009e6
    );
  blk00000900 : XORCY
    port map (
      CI => sig000009e4,
      LI => sig000009e5,
      O => sig00000891
    );
  blk00000901 : LUT2
    generic map(
      INIT => X"9"
    )
    port map (
      I0 => sig000007ec,
      I1 => sig0000082a,
      O => sig000009e7
    );
  blk00000902 : MUXCY
    port map (
      CI => sig000009e6,
      DI => sig000007ec,
      S => sig000009e7,
      O => sig000009e8
    );
  blk00000903 : XORCY
    port map (
      CI => sig000009e6,
      LI => sig000009e7,
      O => sig00000890
    );
  blk00000904 : LUT2
    generic map(
      INIT => X"9"
    )
    port map (
      I0 => sig000007eb,
      I1 => sig00000829,
      O => sig000009e9
    );
  blk00000905 : MUXCY
    port map (
      CI => sig000009e8,
      DI => sig000007eb,
      S => sig000009e9,
      O => sig000009ea
    );
  blk00000906 : XORCY
    port map (
      CI => sig000009e8,
      LI => sig000009e9,
      O => sig0000088f
    );
  blk00000907 : LUT2
    generic map(
      INIT => X"9"
    )
    port map (
      I0 => sig000007ea,
      I1 => sig00000828,
      O => sig000009eb
    );
  blk00000908 : MUXCY
    port map (
      CI => sig000009ea,
      DI => sig000007ea,
      S => sig000009eb,
      O => sig000009ec
    );
  blk00000909 : XORCY
    port map (
      CI => sig000009ea,
      LI => sig000009eb,
      O => sig0000088e
    );
  blk0000090a : LUT2
    generic map(
      INIT => X"9"
    )
    port map (
      I0 => sig000007e9,
      I1 => sig00000827,
      O => sig000009ed
    );
  blk0000090b : MUXCY
    port map (
      CI => sig000009ec,
      DI => sig000007e9,
      S => sig000009ed,
      O => sig000009ee
    );
  blk0000090c : XORCY
    port map (
      CI => sig000009ec,
      LI => sig000009ed,
      O => sig0000088d
    );
  blk0000090d : LUT2
    generic map(
      INIT => X"9"
    )
    port map (
      I0 => sig000007e8,
      I1 => sig00000826,
      O => sig000009ef
    );
  blk0000090e : MUXCY
    port map (
      CI => sig000009ee,
      DI => sig000007e8,
      S => sig000009ef,
      O => sig000009f0
    );
  blk0000090f : XORCY
    port map (
      CI => sig000009ee,
      LI => sig000009ef,
      O => sig0000088c
    );
  blk00000910 : LUT2
    generic map(
      INIT => X"9"
    )
    port map (
      I0 => sig000007e7,
      I1 => sig00000825,
      O => sig000009f1
    );
  blk00000911 : MUXCY
    port map (
      CI => sig000009f0,
      DI => sig000007e7,
      S => sig000009f1,
      O => sig000009f2
    );
  blk00000912 : XORCY
    port map (
      CI => sig000009f0,
      LI => sig000009f1,
      O => sig0000088b
    );
  blk00000913 : LUT2
    generic map(
      INIT => X"9"
    )
    port map (
      I0 => sig000007e6,
      I1 => sig00000824,
      O => sig000009f3
    );
  blk00000914 : MUXCY
    port map (
      CI => sig000009f2,
      DI => sig000007e6,
      S => sig00000ef2,
      O => sig000009f4
    );
  blk00000915 : XORCY
    port map (
      CI => sig000009f2,
      LI => sig00000ef2,
      O => sig0000088a
    );
  blk00000916 : XORCY
    port map (
      CI => sig000009f4,
      LI => sig000009f3,
      O => sig00000889
    );
  blk00000917 : DSP48E
    generic map(
      ACASCREG => 2,
      ALUMODEREG => 0,
      AREG => 2,
      AUTORESET_PATTERN_DETECT => FALSE,
      AUTORESET_PATTERN_DETECT_OPTINV => "MATCH",
      A_INPUT => "DIRECT",
      BCASCREG => 2,
      BREG => 2,
      B_INPUT => "DIRECT",
      CARRYINREG => 0,
      CARRYINSELREG => 0,
      CREG => 1,
      MASK => X"000000000000",
      MREG => 1,
      MULTCARRYINREG => 0,
      OPMODEREG => 0,
      PATTERN => X"000000000000",
      PREG => 1,
      SEL_MASK => "MASK",
      SEL_PATTERN => "PATTERN",
      SEL_ROUNDING_MASK => "SEL_MASK",
      SIM_MODE => "SAFE",
      USE_MULT => "MULT_S",
      USE_PATTERN_DETECT => "NO_PATDET",
      USE_SIMD => "ONE48"
    )
    port map (
      CARRYIN => sig000008b6,
      CEA1 => ce,
      CEA2 => ce,
      CEB1 => ce,
      CEB2 => ce,
      CEC => ce,
      CECTRL => sig000008b6,
      CEP => ce,
      CEM => ce,
      CECARRYIN => sig000008b6,
      CEMULTCARRYIN => sig000008b6,
      CLK => clk,
      RSTA => sig000008b6,
      RSTB => sig000008b6,
      RSTC => sig000008b6,
      RSTCTRL => sig000008b6,
      RSTP => sig000008b6,
      RSTM => sig000008b6,
      RSTALLCARRYIN => sig000008b6,
      CEALUMODE => sig000008b6,
      RSTALUMODE => sig000008b6,
      PATTERNBDETECT => NLW_blk00000917_PATTERNBDETECT_UNCONNECTED,
      PATTERNDETECT => NLW_blk00000917_PATTERNDETECT_UNCONNECTED,
      OVERFLOW => NLW_blk00000917_OVERFLOW_UNCONNECTED,
      UNDERFLOW => NLW_blk00000917_UNDERFLOW_UNCONNECTED,
      CARRYCASCIN => sig000008b6,
      CARRYCASCOUT => NLW_blk00000917_CARRYCASCOUT_UNCONNECTED,
      MULTSIGNIN => sig000008b6,
      MULTSIGNOUT => NLW_blk00000917_MULTSIGNOUT_UNCONNECTED,
      A(29) => sig000008b6,
      A(28) => sig000008b6,
      A(27) => sig000008b6,
      A(26) => sig000008b6,
      A(25) => sig000008b6,
      A(24) => sig00000819,
      A(23) => sig00000819,
      A(22) => sig00000819,
      A(21) => sig00000819,
      A(20) => sig00000819,
      A(19) => sig00000819,
      A(18) => sig00000819,
      A(17) => sig00000819,
      A(16) => sig00000819,
      A(15) => sig00000819,
      A(14) => sig00000819,
      A(13) => sig00000819,
      A(12) => sig00000819,
      A(11) => sig0000081a,
      A(10) => sig0000081b,
      A(9) => sig0000081c,
      A(8) => sig0000081d,
      A(7) => sig0000081e,
      A(6) => sig0000081f,
      A(5) => sig00000820,
      A(4) => sig00000821,
      A(3) => sig00000822,
      A(2) => sig00000823,
      A(1) => sig000008b6,
      A(0) => sig000008b6,
      PCIN(47) => sig000008b6,
      PCIN(46) => sig000008b6,
      PCIN(45) => sig000008b6,
      PCIN(44) => sig000008b6,
      PCIN(43) => sig000008b6,
      PCIN(42) => sig000008b6,
      PCIN(41) => sig000008b6,
      PCIN(40) => sig000008b6,
      PCIN(39) => sig000008b6,
      PCIN(38) => sig000008b6,
      PCIN(37) => sig000008b6,
      PCIN(36) => sig000008b6,
      PCIN(35) => sig000008b6,
      PCIN(34) => sig000008b6,
      PCIN(33) => sig000008b6,
      PCIN(32) => sig000008b6,
      PCIN(31) => sig000008b6,
      PCIN(30) => sig000008b6,
      PCIN(29) => sig000008b6,
      PCIN(28) => sig000008b6,
      PCIN(27) => sig000008b6,
      PCIN(26) => sig000008b6,
      PCIN(25) => sig000008b6,
      PCIN(24) => sig000008b6,
      PCIN(23) => sig000008b6,
      PCIN(22) => sig000008b6,
      PCIN(21) => sig000008b6,
      PCIN(20) => sig000008b6,
      PCIN(19) => sig000008b6,
      PCIN(18) => sig000008b6,
      PCIN(17) => sig000008b6,
      PCIN(16) => sig000008b6,
      PCIN(15) => sig000008b6,
      PCIN(14) => sig000008b6,
      PCIN(13) => sig000008b6,
      PCIN(12) => sig000008b6,
      PCIN(11) => sig000008b6,
      PCIN(10) => sig000008b6,
      PCIN(9) => sig000008b6,
      PCIN(8) => sig000008b6,
      PCIN(7) => sig000008b6,
      PCIN(6) => sig000008b6,
      PCIN(5) => sig000008b6,
      PCIN(4) => sig000008b6,
      PCIN(3) => sig000008b6,
      PCIN(2) => sig000008b6,
      PCIN(1) => sig000008b6,
      PCIN(0) => sig000008b6,
      B(17) => sig0000080a,
      B(16) => sig0000080a,
      B(15) => sig0000080a,
      B(14) => sig0000080a,
      B(13) => sig0000080b,
      B(12) => sig0000080c,
      B(11) => sig0000080d,
      B(10) => sig0000080e,
      B(9) => sig0000080f,
      B(8) => sig00000810,
      B(7) => sig00000811,
      B(6) => sig00000812,
      B(5) => sig00000813,
      B(4) => sig00000814,
      B(3) => sig00000815,
      B(2) => sig00000816,
      B(1) => sig00000817,
      B(0) => sig00000818,
      C(47) => sig00000832,
      C(46) => sig00000832,
      C(45) => sig00000832,
      C(44) => sig00000832,
      C(43) => sig00000832,
      C(42) => sig00000832,
      C(41) => sig00000832,
      C(40) => sig00000832,
      C(39) => sig00000832,
      C(38) => sig00000832,
      C(37) => sig00000832,
      C(36) => sig00000832,
      C(35) => sig00000832,
      C(34) => sig00000832,
      C(33) => sig00000832,
      C(32) => sig00000832,
      C(31) => sig00000832,
      C(30) => sig00000832,
      C(29) => sig00000832,
      C(28) => sig00000832,
      C(27) => sig00000832,
      C(26) => sig00000833,
      C(25) => sig00000834,
      C(24) => sig00000835,
      C(23) => sig00000836,
      C(22) => sig00000837,
      C(21) => sig00000838,
      C(20) => sig00000839,
      C(19) => sig0000083a,
      C(18) => sig0000083b,
      C(17) => sig0000083c,
      C(16) => sig0000083d,
      C(15) => sig0000083e,
      C(14) => sig0000083f,
      C(13) => sig00000840,
      C(12) => sig00000841,
      C(11) => sig00000842,
      C(10) => sig00000843,
      C(9) => sig00000844,
      C(8) => sig00000845,
      C(7) => sig00000846,
      C(6) => sig00000847,
      C(5) => sig00000848,
      C(4) => sig00000849,
      C(3) => sig0000084a,
      C(2) => sig0000084b,
      C(1) => sig0000084c,
      C(0) => sig0000084d,
      CARRYINSEL(2) => sig000008b6,
      CARRYINSEL(1) => sig000008b6,
      CARRYINSEL(0) => sig000008b6,
      OPMODE(6) => sig000008b6,
      OPMODE(5) => sig000006d1,
      OPMODE(4) => sig000006d1,
      OPMODE(3) => sig000008b6,
      OPMODE(2) => sig000006d1,
      OPMODE(1) => sig000008b6,
      OPMODE(0) => sig000006d1,
      BCIN(17) => sig000008b6,
      BCIN(16) => sig000008b6,
      BCIN(15) => sig000008b6,
      BCIN(14) => sig000008b6,
      BCIN(13) => sig000008b6,
      BCIN(12) => sig000008b6,
      BCIN(11) => sig000008b6,
      BCIN(10) => sig000008b6,
      BCIN(9) => sig000008b6,
      BCIN(8) => sig000008b6,
      BCIN(7) => sig000008b6,
      BCIN(6) => sig000008b6,
      BCIN(5) => sig000008b6,
      BCIN(4) => sig000008b6,
      BCIN(3) => sig000008b6,
      BCIN(2) => sig000008b6,
      BCIN(1) => sig000008b6,
      BCIN(0) => sig000008b6,
      ALUMODE(3) => sig000008b6,
      ALUMODE(2) => sig000008b6,
      ALUMODE(1) => sig000006d1,
      ALUMODE(0) => sig000006d1,
      PCOUT(47) => NLW_blk00000917_PCOUT_47_UNCONNECTED,
      PCOUT(46) => NLW_blk00000917_PCOUT_46_UNCONNECTED,
      PCOUT(45) => NLW_blk00000917_PCOUT_45_UNCONNECTED,
      PCOUT(44) => NLW_blk00000917_PCOUT_44_UNCONNECTED,
      PCOUT(43) => NLW_blk00000917_PCOUT_43_UNCONNECTED,
      PCOUT(42) => NLW_blk00000917_PCOUT_42_UNCONNECTED,
      PCOUT(41) => NLW_blk00000917_PCOUT_41_UNCONNECTED,
      PCOUT(40) => NLW_blk00000917_PCOUT_40_UNCONNECTED,
      PCOUT(39) => NLW_blk00000917_PCOUT_39_UNCONNECTED,
      PCOUT(38) => NLW_blk00000917_PCOUT_38_UNCONNECTED,
      PCOUT(37) => NLW_blk00000917_PCOUT_37_UNCONNECTED,
      PCOUT(36) => NLW_blk00000917_PCOUT_36_UNCONNECTED,
      PCOUT(35) => NLW_blk00000917_PCOUT_35_UNCONNECTED,
      PCOUT(34) => NLW_blk00000917_PCOUT_34_UNCONNECTED,
      PCOUT(33) => NLW_blk00000917_PCOUT_33_UNCONNECTED,
      PCOUT(32) => NLW_blk00000917_PCOUT_32_UNCONNECTED,
      PCOUT(31) => NLW_blk00000917_PCOUT_31_UNCONNECTED,
      PCOUT(30) => NLW_blk00000917_PCOUT_30_UNCONNECTED,
      PCOUT(29) => NLW_blk00000917_PCOUT_29_UNCONNECTED,
      PCOUT(28) => NLW_blk00000917_PCOUT_28_UNCONNECTED,
      PCOUT(27) => NLW_blk00000917_PCOUT_27_UNCONNECTED,
      PCOUT(26) => NLW_blk00000917_PCOUT_26_UNCONNECTED,
      PCOUT(25) => NLW_blk00000917_PCOUT_25_UNCONNECTED,
      PCOUT(24) => NLW_blk00000917_PCOUT_24_UNCONNECTED,
      PCOUT(23) => NLW_blk00000917_PCOUT_23_UNCONNECTED,
      PCOUT(22) => NLW_blk00000917_PCOUT_22_UNCONNECTED,
      PCOUT(21) => NLW_blk00000917_PCOUT_21_UNCONNECTED,
      PCOUT(20) => NLW_blk00000917_PCOUT_20_UNCONNECTED,
      PCOUT(19) => NLW_blk00000917_PCOUT_19_UNCONNECTED,
      PCOUT(18) => NLW_blk00000917_PCOUT_18_UNCONNECTED,
      PCOUT(17) => NLW_blk00000917_PCOUT_17_UNCONNECTED,
      PCOUT(16) => NLW_blk00000917_PCOUT_16_UNCONNECTED,
      PCOUT(15) => NLW_blk00000917_PCOUT_15_UNCONNECTED,
      PCOUT(14) => NLW_blk00000917_PCOUT_14_UNCONNECTED,
      PCOUT(13) => NLW_blk00000917_PCOUT_13_UNCONNECTED,
      PCOUT(12) => NLW_blk00000917_PCOUT_12_UNCONNECTED,
      PCOUT(11) => NLW_blk00000917_PCOUT_11_UNCONNECTED,
      PCOUT(10) => NLW_blk00000917_PCOUT_10_UNCONNECTED,
      PCOUT(9) => NLW_blk00000917_PCOUT_9_UNCONNECTED,
      PCOUT(8) => NLW_blk00000917_PCOUT_8_UNCONNECTED,
      PCOUT(7) => NLW_blk00000917_PCOUT_7_UNCONNECTED,
      PCOUT(6) => NLW_blk00000917_PCOUT_6_UNCONNECTED,
      PCOUT(5) => NLW_blk00000917_PCOUT_5_UNCONNECTED,
      PCOUT(4) => NLW_blk00000917_PCOUT_4_UNCONNECTED,
      PCOUT(3) => NLW_blk00000917_PCOUT_3_UNCONNECTED,
      PCOUT(2) => NLW_blk00000917_PCOUT_2_UNCONNECTED,
      PCOUT(1) => NLW_blk00000917_PCOUT_1_UNCONNECTED,
      PCOUT(0) => NLW_blk00000917_PCOUT_0_UNCONNECTED,
      P(47) => NLW_blk00000917_P_47_UNCONNECTED,
      P(46) => NLW_blk00000917_P_46_UNCONNECTED,
      P(45) => NLW_blk00000917_P_45_UNCONNECTED,
      P(44) => NLW_blk00000917_P_44_UNCONNECTED,
      P(43) => NLW_blk00000917_P_43_UNCONNECTED,
      P(42) => sig000008f9,
      P(41) => sig000008f8,
      P(40) => sig000008f7,
      P(39) => sig000008f6,
      P(38) => sig000008f5,
      P(37) => sig000008f4,
      P(36) => sig000008f3,
      P(35) => sig000008f2,
      P(34) => sig000008f1,
      P(33) => sig000008f0,
      P(32) => sig000008ef,
      P(31) => sig000008ee,
      P(30) => sig000008ed,
      P(29) => sig000008ec,
      P(28) => sig000008eb,
      P(27) => sig000008ea,
      P(26) => sig000008e9,
      P(25) => sig000008e8,
      P(24) => sig000008e7,
      P(23) => sig000008e6,
      P(22) => sig000008e5,
      P(21) => sig000008e4,
      P(20) => sig000008e3,
      P(19) => sig000008e2,
      P(18) => sig000008e1,
      P(17) => sig000008e0,
      P(16) => sig000008df,
      P(15) => sig000008de,
      P(14) => sig000008dd,
      P(13) => sig000008dc,
      P(12) => sig000008db,
      P(11) => sig000008da,
      P(10) => sig000008d9,
      P(9) => sig000008d8,
      P(8) => sig000008d7,
      P(7) => sig000008d6,
      P(6) => sig000008d5,
      P(5) => sig000008d4,
      P(4) => sig000008d3,
      P(3) => sig000008d2,
      P(2) => sig000008d1,
      P(1) => sig000008d0,
      P(0) => sig000008cf,
      BCOUT(17) => NLW_blk00000917_BCOUT_17_UNCONNECTED,
      BCOUT(16) => NLW_blk00000917_BCOUT_16_UNCONNECTED,
      BCOUT(15) => NLW_blk00000917_BCOUT_15_UNCONNECTED,
      BCOUT(14) => NLW_blk00000917_BCOUT_14_UNCONNECTED,
      BCOUT(13) => NLW_blk00000917_BCOUT_13_UNCONNECTED,
      BCOUT(12) => NLW_blk00000917_BCOUT_12_UNCONNECTED,
      BCOUT(11) => NLW_blk00000917_BCOUT_11_UNCONNECTED,
      BCOUT(10) => NLW_blk00000917_BCOUT_10_UNCONNECTED,
      BCOUT(9) => NLW_blk00000917_BCOUT_9_UNCONNECTED,
      BCOUT(8) => NLW_blk00000917_BCOUT_8_UNCONNECTED,
      BCOUT(7) => NLW_blk00000917_BCOUT_7_UNCONNECTED,
      BCOUT(6) => NLW_blk00000917_BCOUT_6_UNCONNECTED,
      BCOUT(5) => NLW_blk00000917_BCOUT_5_UNCONNECTED,
      BCOUT(4) => NLW_blk00000917_BCOUT_4_UNCONNECTED,
      BCOUT(3) => NLW_blk00000917_BCOUT_3_UNCONNECTED,
      BCOUT(2) => NLW_blk00000917_BCOUT_2_UNCONNECTED,
      BCOUT(1) => NLW_blk00000917_BCOUT_1_UNCONNECTED,
      BCOUT(0) => NLW_blk00000917_BCOUT_0_UNCONNECTED,
      ACIN(29) => sig000008b6,
      ACIN(28) => sig000008b6,
      ACIN(27) => sig000008b6,
      ACIN(26) => sig000008b6,
      ACIN(25) => sig000008b6,
      ACIN(24) => sig000008b6,
      ACIN(23) => sig000008b6,
      ACIN(22) => sig000008b6,
      ACIN(21) => sig000008b6,
      ACIN(20) => sig000008b6,
      ACIN(19) => sig000008b6,
      ACIN(18) => sig000008b6,
      ACIN(17) => sig000008b6,
      ACIN(16) => sig000008b6,
      ACIN(15) => sig000008b6,
      ACIN(14) => sig000008b6,
      ACIN(13) => sig000008b6,
      ACIN(12) => sig000008b6,
      ACIN(11) => sig000008b6,
      ACIN(10) => sig000008b6,
      ACIN(9) => sig000008b6,
      ACIN(8) => sig000008b6,
      ACIN(7) => sig000008b6,
      ACIN(6) => sig000008b6,
      ACIN(5) => sig000008b6,
      ACIN(4) => sig000008b6,
      ACIN(3) => sig000008b6,
      ACIN(2) => sig000008b6,
      ACIN(1) => sig000008b6,
      ACIN(0) => sig000008b6,
      ACOUT(29) => NLW_blk00000917_ACOUT_29_UNCONNECTED,
      ACOUT(28) => NLW_blk00000917_ACOUT_28_UNCONNECTED,
      ACOUT(27) => NLW_blk00000917_ACOUT_27_UNCONNECTED,
      ACOUT(26) => NLW_blk00000917_ACOUT_26_UNCONNECTED,
      ACOUT(25) => NLW_blk00000917_ACOUT_25_UNCONNECTED,
      ACOUT(24) => NLW_blk00000917_ACOUT_24_UNCONNECTED,
      ACOUT(23) => NLW_blk00000917_ACOUT_23_UNCONNECTED,
      ACOUT(22) => NLW_blk00000917_ACOUT_22_UNCONNECTED,
      ACOUT(21) => NLW_blk00000917_ACOUT_21_UNCONNECTED,
      ACOUT(20) => NLW_blk00000917_ACOUT_20_UNCONNECTED,
      ACOUT(19) => NLW_blk00000917_ACOUT_19_UNCONNECTED,
      ACOUT(18) => NLW_blk00000917_ACOUT_18_UNCONNECTED,
      ACOUT(17) => NLW_blk00000917_ACOUT_17_UNCONNECTED,
      ACOUT(16) => NLW_blk00000917_ACOUT_16_UNCONNECTED,
      ACOUT(15) => NLW_blk00000917_ACOUT_15_UNCONNECTED,
      ACOUT(14) => NLW_blk00000917_ACOUT_14_UNCONNECTED,
      ACOUT(13) => NLW_blk00000917_ACOUT_13_UNCONNECTED,
      ACOUT(12) => NLW_blk00000917_ACOUT_12_UNCONNECTED,
      ACOUT(11) => NLW_blk00000917_ACOUT_11_UNCONNECTED,
      ACOUT(10) => NLW_blk00000917_ACOUT_10_UNCONNECTED,
      ACOUT(9) => NLW_blk00000917_ACOUT_9_UNCONNECTED,
      ACOUT(8) => NLW_blk00000917_ACOUT_8_UNCONNECTED,
      ACOUT(7) => NLW_blk00000917_ACOUT_7_UNCONNECTED,
      ACOUT(6) => NLW_blk00000917_ACOUT_6_UNCONNECTED,
      ACOUT(5) => NLW_blk00000917_ACOUT_5_UNCONNECTED,
      ACOUT(4) => NLW_blk00000917_ACOUT_4_UNCONNECTED,
      ACOUT(3) => NLW_blk00000917_ACOUT_3_UNCONNECTED,
      ACOUT(2) => NLW_blk00000917_ACOUT_2_UNCONNECTED,
      ACOUT(1) => NLW_blk00000917_ACOUT_1_UNCONNECTED,
      ACOUT(0) => NLW_blk00000917_ACOUT_0_UNCONNECTED,
      CARRYOUT(3) => NLW_blk00000917_CARRYOUT_3_UNCONNECTED,
      CARRYOUT(2) => NLW_blk00000917_CARRYOUT_2_UNCONNECTED,
      CARRYOUT(1) => NLW_blk00000917_CARRYOUT_1_UNCONNECTED,
      CARRYOUT(0) => NLW_blk00000917_CARRYOUT_0_UNCONNECTED
    );
  blk00000918 : DSP48E
    generic map(
      ACASCREG => 2,
      ALUMODEREG => 0,
      AREG => 2,
      AUTORESET_PATTERN_DETECT => FALSE,
      AUTORESET_PATTERN_DETECT_OPTINV => "MATCH",
      A_INPUT => "DIRECT",
      BCASCREG => 1,
      BREG => 1,
      B_INPUT => "DIRECT",
      CARRYINREG => 0,
      CARRYINSELREG => 0,
      CREG => 0,
      MASK => X"000000000000",
      MREG => 1,
      MULTCARRYINREG => 0,
      OPMODEREG => 0,
      PATTERN => X"000000000000",
      PREG => 1,
      SEL_MASK => "MASK",
      SEL_PATTERN => "PATTERN",
      SEL_ROUNDING_MASK => "SEL_MASK",
      SIM_MODE => "SAFE",
      USE_MULT => "MULT_S",
      USE_PATTERN_DETECT => "NO_PATDET",
      USE_SIMD => "ONE48"
    )
    port map (
      CARRYIN => sig000008b6,
      CEA1 => ce,
      CEA2 => ce,
      CEB1 => sig000008b6,
      CEB2 => ce,
      CEC => sig000008b6,
      CECTRL => sig000008b6,
      CEP => ce,
      CEM => ce,
      CECARRYIN => sig000008b6,
      CEMULTCARRYIN => sig000008b6,
      CLK => clk,
      RSTA => sig000008b6,
      RSTB => sig000008b6,
      RSTC => sig000008b6,
      RSTCTRL => sig000008b6,
      RSTP => sig000008b6,
      RSTM => sig000008b6,
      RSTALLCARRYIN => sig000008b6,
      CEALUMODE => sig000008b6,
      RSTALUMODE => sig000008b6,
      PATTERNBDETECT => NLW_blk00000918_PATTERNBDETECT_UNCONNECTED,
      PATTERNDETECT => NLW_blk00000918_PATTERNDETECT_UNCONNECTED,
      OVERFLOW => NLW_blk00000918_OVERFLOW_UNCONNECTED,
      UNDERFLOW => NLW_blk00000918_UNDERFLOW_UNCONNECTED,
      CARRYCASCIN => sig000008b6,
      CARRYCASCOUT => NLW_blk00000918_CARRYCASCOUT_UNCONNECTED,
      MULTSIGNIN => sig000008b6,
      MULTSIGNOUT => NLW_blk00000918_MULTSIGNOUT_UNCONNECTED,
      A(29) => sig000008b6,
      A(28) => sig000008b6,
      A(27) => sig000008b6,
      A(26) => sig000008b6,
      A(25) => sig000008b6,
      A(24) => sig00000824,
      A(23) => sig00000824,
      A(22) => sig00000824,
      A(21) => sig00000824,
      A(20) => sig00000824,
      A(19) => sig00000824,
      A(18) => sig00000824,
      A(17) => sig00000824,
      A(16) => sig00000824,
      A(15) => sig00000824,
      A(14) => sig00000824,
      A(13) => sig00000824,
      A(12) => sig00000825,
      A(11) => sig00000826,
      A(10) => sig00000827,
      A(9) => sig00000828,
      A(8) => sig00000829,
      A(7) => sig0000082a,
      A(6) => sig0000082b,
      A(5) => sig0000082c,
      A(4) => sig0000082d,
      A(3) => sig0000082e,
      A(2) => sig0000082f,
      A(1) => sig00000830,
      A(0) => sig00000831,
      PCIN(47) => sig000008b6,
      PCIN(46) => sig000008b6,
      PCIN(45) => sig000008b6,
      PCIN(44) => sig000008b6,
      PCIN(43) => sig000008b6,
      PCIN(42) => sig000008b6,
      PCIN(41) => sig000008b6,
      PCIN(40) => sig000008b6,
      PCIN(39) => sig000008b6,
      PCIN(38) => sig000008b6,
      PCIN(37) => sig000008b6,
      PCIN(36) => sig000008b6,
      PCIN(35) => sig000008b6,
      PCIN(34) => sig000008b6,
      PCIN(33) => sig000008b6,
      PCIN(32) => sig000008b6,
      PCIN(31) => sig000008b6,
      PCIN(30) => sig000008b6,
      PCIN(29) => sig000008b6,
      PCIN(28) => sig000008b6,
      PCIN(27) => sig000008b6,
      PCIN(26) => sig000008b6,
      PCIN(25) => sig000008b6,
      PCIN(24) => sig000008b6,
      PCIN(23) => sig000008b6,
      PCIN(22) => sig000008b6,
      PCIN(21) => sig000008b6,
      PCIN(20) => sig000008b6,
      PCIN(19) => sig000008b6,
      PCIN(18) => sig000008b6,
      PCIN(17) => sig000008b6,
      PCIN(16) => sig000008b6,
      PCIN(15) => sig000008b6,
      PCIN(14) => sig000008b6,
      PCIN(13) => sig000008b6,
      PCIN(12) => sig000008b6,
      PCIN(11) => sig000008b6,
      PCIN(10) => sig000008b6,
      PCIN(9) => sig000008b6,
      PCIN(8) => sig000008b6,
      PCIN(7) => sig000008b6,
      PCIN(6) => sig000008b6,
      PCIN(5) => sig000008b6,
      PCIN(4) => sig000008b6,
      PCIN(3) => sig000008b6,
      PCIN(2) => sig000008b6,
      PCIN(1) => sig000008b6,
      PCIN(0) => sig000008b6,
      B(17) => sig00000867,
      B(16) => sig00000867,
      B(15) => sig00000867,
      B(14) => sig00000867,
      B(13) => sig00000867,
      B(12) => sig00000868,
      B(11) => sig00000869,
      B(10) => sig0000086a,
      B(9) => sig0000086b,
      B(8) => sig0000086c,
      B(7) => sig0000086d,
      B(6) => sig0000086e,
      B(5) => sig0000086f,
      B(4) => sig00000870,
      B(3) => sig00000871,
      B(2) => sig00000872,
      B(1) => sig000008b6,
      B(0) => sig000008b6,
      C(47) => sig000008b6,
      C(46) => sig000008b6,
      C(45) => sig000008b6,
      C(44) => sig000008b6,
      C(43) => sig000008b6,
      C(42) => sig000008b6,
      C(41) => sig000008b6,
      C(40) => sig000008b6,
      C(39) => sig000008b6,
      C(38) => sig000008b6,
      C(37) => sig000008b6,
      C(36) => sig000008b6,
      C(35) => sig000008b6,
      C(34) => sig000008b6,
      C(33) => sig000008b6,
      C(32) => sig000008b6,
      C(31) => sig000008b6,
      C(30) => sig000008b6,
      C(29) => sig000008b6,
      C(28) => sig000008b6,
      C(27) => sig000008b6,
      C(26) => sig000008b6,
      C(25) => sig000008b6,
      C(24) => sig000008b6,
      C(23) => sig000008b6,
      C(22) => sig000008b6,
      C(21) => sig000008b6,
      C(20) => sig000008b6,
      C(19) => sig000008b6,
      C(18) => sig000008b6,
      C(17) => sig000008b6,
      C(16) => sig000008b6,
      C(15) => sig000008b6,
      C(14) => sig000008b6,
      C(13) => sig000008b6,
      C(12) => sig000008b6,
      C(11) => sig000008b6,
      C(10) => sig000008b6,
      C(9) => sig000008b6,
      C(8) => sig000008b6,
      C(7) => sig000008b6,
      C(6) => sig000008b6,
      C(5) => sig000008b6,
      C(4) => sig000006d1,
      C(3) => sig000006d1,
      C(2) => sig000006d1,
      C(1) => sig000006d1,
      C(0) => sig000006d1,
      CARRYINSEL(2) => sig000008b6,
      CARRYINSEL(1) => sig000008b6,
      CARRYINSEL(0) => sig000008b6,
      OPMODE(6) => sig000008b6,
      OPMODE(5) => sig000006d1,
      OPMODE(4) => sig000006d1,
      OPMODE(3) => sig000008b6,
      OPMODE(2) => sig000006d1,
      OPMODE(1) => sig000008b6,
      OPMODE(0) => sig000006d1,
      BCIN(17) => sig000008b6,
      BCIN(16) => sig000008b6,
      BCIN(15) => sig000008b6,
      BCIN(14) => sig000008b6,
      BCIN(13) => sig000008b6,
      BCIN(12) => sig000008b6,
      BCIN(11) => sig000008b6,
      BCIN(10) => sig000008b6,
      BCIN(9) => sig000008b6,
      BCIN(8) => sig000008b6,
      BCIN(7) => sig000008b6,
      BCIN(6) => sig000008b6,
      BCIN(5) => sig000008b6,
      BCIN(4) => sig000008b6,
      BCIN(3) => sig000008b6,
      BCIN(2) => sig000008b6,
      BCIN(1) => sig000008b6,
      BCIN(0) => sig000008b6,
      ALUMODE(3) => sig000008b6,
      ALUMODE(2) => sig000008b6,
      ALUMODE(1) => sig000008b6,
      ALUMODE(0) => sig000008b6,
      PCOUT(47) => NLW_blk00000918_PCOUT_47_UNCONNECTED,
      PCOUT(46) => NLW_blk00000918_PCOUT_46_UNCONNECTED,
      PCOUT(45) => NLW_blk00000918_PCOUT_45_UNCONNECTED,
      PCOUT(44) => NLW_blk00000918_PCOUT_44_UNCONNECTED,
      PCOUT(43) => NLW_blk00000918_PCOUT_43_UNCONNECTED,
      PCOUT(42) => NLW_blk00000918_PCOUT_42_UNCONNECTED,
      PCOUT(41) => NLW_blk00000918_PCOUT_41_UNCONNECTED,
      PCOUT(40) => NLW_blk00000918_PCOUT_40_UNCONNECTED,
      PCOUT(39) => NLW_blk00000918_PCOUT_39_UNCONNECTED,
      PCOUT(38) => NLW_blk00000918_PCOUT_38_UNCONNECTED,
      PCOUT(37) => NLW_blk00000918_PCOUT_37_UNCONNECTED,
      PCOUT(36) => NLW_blk00000918_PCOUT_36_UNCONNECTED,
      PCOUT(35) => NLW_blk00000918_PCOUT_35_UNCONNECTED,
      PCOUT(34) => NLW_blk00000918_PCOUT_34_UNCONNECTED,
      PCOUT(33) => NLW_blk00000918_PCOUT_33_UNCONNECTED,
      PCOUT(32) => NLW_blk00000918_PCOUT_32_UNCONNECTED,
      PCOUT(31) => NLW_blk00000918_PCOUT_31_UNCONNECTED,
      PCOUT(30) => NLW_blk00000918_PCOUT_30_UNCONNECTED,
      PCOUT(29) => NLW_blk00000918_PCOUT_29_UNCONNECTED,
      PCOUT(28) => NLW_blk00000918_PCOUT_28_UNCONNECTED,
      PCOUT(27) => NLW_blk00000918_PCOUT_27_UNCONNECTED,
      PCOUT(26) => NLW_blk00000918_PCOUT_26_UNCONNECTED,
      PCOUT(25) => NLW_blk00000918_PCOUT_25_UNCONNECTED,
      PCOUT(24) => NLW_blk00000918_PCOUT_24_UNCONNECTED,
      PCOUT(23) => NLW_blk00000918_PCOUT_23_UNCONNECTED,
      PCOUT(22) => NLW_blk00000918_PCOUT_22_UNCONNECTED,
      PCOUT(21) => NLW_blk00000918_PCOUT_21_UNCONNECTED,
      PCOUT(20) => NLW_blk00000918_PCOUT_20_UNCONNECTED,
      PCOUT(19) => NLW_blk00000918_PCOUT_19_UNCONNECTED,
      PCOUT(18) => NLW_blk00000918_PCOUT_18_UNCONNECTED,
      PCOUT(17) => NLW_blk00000918_PCOUT_17_UNCONNECTED,
      PCOUT(16) => NLW_blk00000918_PCOUT_16_UNCONNECTED,
      PCOUT(15) => NLW_blk00000918_PCOUT_15_UNCONNECTED,
      PCOUT(14) => NLW_blk00000918_PCOUT_14_UNCONNECTED,
      PCOUT(13) => NLW_blk00000918_PCOUT_13_UNCONNECTED,
      PCOUT(12) => NLW_blk00000918_PCOUT_12_UNCONNECTED,
      PCOUT(11) => NLW_blk00000918_PCOUT_11_UNCONNECTED,
      PCOUT(10) => NLW_blk00000918_PCOUT_10_UNCONNECTED,
      PCOUT(9) => NLW_blk00000918_PCOUT_9_UNCONNECTED,
      PCOUT(8) => NLW_blk00000918_PCOUT_8_UNCONNECTED,
      PCOUT(7) => NLW_blk00000918_PCOUT_7_UNCONNECTED,
      PCOUT(6) => NLW_blk00000918_PCOUT_6_UNCONNECTED,
      PCOUT(5) => NLW_blk00000918_PCOUT_5_UNCONNECTED,
      PCOUT(4) => NLW_blk00000918_PCOUT_4_UNCONNECTED,
      PCOUT(3) => NLW_blk00000918_PCOUT_3_UNCONNECTED,
      PCOUT(2) => NLW_blk00000918_PCOUT_2_UNCONNECTED,
      PCOUT(1) => NLW_blk00000918_PCOUT_1_UNCONNECTED,
      PCOUT(0) => NLW_blk00000918_PCOUT_0_UNCONNECTED,
      P(47) => NLW_blk00000918_P_47_UNCONNECTED,
      P(46) => NLW_blk00000918_P_46_UNCONNECTED,
      P(45) => NLW_blk00000918_P_45_UNCONNECTED,
      P(44) => NLW_blk00000918_P_44_UNCONNECTED,
      P(43) => NLW_blk00000918_P_43_UNCONNECTED,
      P(42) => sig0000094f,
      P(41) => sig0000094e,
      P(40) => sig0000094d,
      P(39) => sig0000094c,
      P(38) => sig0000094b,
      P(37) => sig0000094a,
      P(36) => sig00000949,
      P(35) => sig00000948,
      P(34) => sig00000947,
      P(33) => sig00000946,
      P(32) => sig00000945,
      P(31) => sig00000944,
      P(30) => sig00000943,
      P(29) => sig00000942,
      P(28) => sig00000941,
      P(27) => sig00000832,
      P(26) => sig00000833,
      P(25) => sig00000834,
      P(24) => sig00000835,
      P(23) => sig00000836,
      P(22) => sig00000837,
      P(21) => sig00000838,
      P(20) => sig00000839,
      P(19) => sig0000083a,
      P(18) => sig0000083b,
      P(17) => sig0000083c,
      P(16) => sig0000083d,
      P(15) => sig0000083e,
      P(14) => sig0000083f,
      P(13) => sig00000840,
      P(12) => sig00000841,
      P(11) => sig00000842,
      P(10) => sig00000843,
      P(9) => sig00000844,
      P(8) => sig00000845,
      P(7) => sig00000846,
      P(6) => sig00000847,
      P(5) => sig00000848,
      P(4) => sig00000849,
      P(3) => sig0000084a,
      P(2) => sig0000084b,
      P(1) => sig0000084c,
      P(0) => sig0000084d,
      BCOUT(17) => NLW_blk00000918_BCOUT_17_UNCONNECTED,
      BCOUT(16) => NLW_blk00000918_BCOUT_16_UNCONNECTED,
      BCOUT(15) => NLW_blk00000918_BCOUT_15_UNCONNECTED,
      BCOUT(14) => NLW_blk00000918_BCOUT_14_UNCONNECTED,
      BCOUT(13) => NLW_blk00000918_BCOUT_13_UNCONNECTED,
      BCOUT(12) => NLW_blk00000918_BCOUT_12_UNCONNECTED,
      BCOUT(11) => NLW_blk00000918_BCOUT_11_UNCONNECTED,
      BCOUT(10) => NLW_blk00000918_BCOUT_10_UNCONNECTED,
      BCOUT(9) => NLW_blk00000918_BCOUT_9_UNCONNECTED,
      BCOUT(8) => NLW_blk00000918_BCOUT_8_UNCONNECTED,
      BCOUT(7) => NLW_blk00000918_BCOUT_7_UNCONNECTED,
      BCOUT(6) => NLW_blk00000918_BCOUT_6_UNCONNECTED,
      BCOUT(5) => NLW_blk00000918_BCOUT_5_UNCONNECTED,
      BCOUT(4) => NLW_blk00000918_BCOUT_4_UNCONNECTED,
      BCOUT(3) => NLW_blk00000918_BCOUT_3_UNCONNECTED,
      BCOUT(2) => NLW_blk00000918_BCOUT_2_UNCONNECTED,
      BCOUT(1) => NLW_blk00000918_BCOUT_1_UNCONNECTED,
      BCOUT(0) => NLW_blk00000918_BCOUT_0_UNCONNECTED,
      ACIN(29) => sig000008b6,
      ACIN(28) => sig000008b6,
      ACIN(27) => sig000008b6,
      ACIN(26) => sig000008b6,
      ACIN(25) => sig000008b6,
      ACIN(24) => sig000008b6,
      ACIN(23) => sig000008b6,
      ACIN(22) => sig000008b6,
      ACIN(21) => sig000008b6,
      ACIN(20) => sig000008b6,
      ACIN(19) => sig000008b6,
      ACIN(18) => sig000008b6,
      ACIN(17) => sig000008b6,
      ACIN(16) => sig000008b6,
      ACIN(15) => sig000008b6,
      ACIN(14) => sig000008b6,
      ACIN(13) => sig000008b6,
      ACIN(12) => sig000008b6,
      ACIN(11) => sig000008b6,
      ACIN(10) => sig000008b6,
      ACIN(9) => sig000008b6,
      ACIN(8) => sig000008b6,
      ACIN(7) => sig000008b6,
      ACIN(6) => sig000008b6,
      ACIN(5) => sig000008b6,
      ACIN(4) => sig000008b6,
      ACIN(3) => sig000008b6,
      ACIN(2) => sig000008b6,
      ACIN(1) => sig000008b6,
      ACIN(0) => sig000008b6,
      ACOUT(29) => NLW_blk00000918_ACOUT_29_UNCONNECTED,
      ACOUT(28) => NLW_blk00000918_ACOUT_28_UNCONNECTED,
      ACOUT(27) => NLW_blk00000918_ACOUT_27_UNCONNECTED,
      ACOUT(26) => NLW_blk00000918_ACOUT_26_UNCONNECTED,
      ACOUT(25) => NLW_blk00000918_ACOUT_25_UNCONNECTED,
      ACOUT(24) => NLW_blk00000918_ACOUT_24_UNCONNECTED,
      ACOUT(23) => NLW_blk00000918_ACOUT_23_UNCONNECTED,
      ACOUT(22) => NLW_blk00000918_ACOUT_22_UNCONNECTED,
      ACOUT(21) => NLW_blk00000918_ACOUT_21_UNCONNECTED,
      ACOUT(20) => NLW_blk00000918_ACOUT_20_UNCONNECTED,
      ACOUT(19) => NLW_blk00000918_ACOUT_19_UNCONNECTED,
      ACOUT(18) => NLW_blk00000918_ACOUT_18_UNCONNECTED,
      ACOUT(17) => NLW_blk00000918_ACOUT_17_UNCONNECTED,
      ACOUT(16) => NLW_blk00000918_ACOUT_16_UNCONNECTED,
      ACOUT(15) => NLW_blk00000918_ACOUT_15_UNCONNECTED,
      ACOUT(14) => NLW_blk00000918_ACOUT_14_UNCONNECTED,
      ACOUT(13) => NLW_blk00000918_ACOUT_13_UNCONNECTED,
      ACOUT(12) => NLW_blk00000918_ACOUT_12_UNCONNECTED,
      ACOUT(11) => NLW_blk00000918_ACOUT_11_UNCONNECTED,
      ACOUT(10) => NLW_blk00000918_ACOUT_10_UNCONNECTED,
      ACOUT(9) => NLW_blk00000918_ACOUT_9_UNCONNECTED,
      ACOUT(8) => NLW_blk00000918_ACOUT_8_UNCONNECTED,
      ACOUT(7) => NLW_blk00000918_ACOUT_7_UNCONNECTED,
      ACOUT(6) => NLW_blk00000918_ACOUT_6_UNCONNECTED,
      ACOUT(5) => NLW_blk00000918_ACOUT_5_UNCONNECTED,
      ACOUT(4) => NLW_blk00000918_ACOUT_4_UNCONNECTED,
      ACOUT(3) => NLW_blk00000918_ACOUT_3_UNCONNECTED,
      ACOUT(2) => NLW_blk00000918_ACOUT_2_UNCONNECTED,
      ACOUT(1) => NLW_blk00000918_ACOUT_1_UNCONNECTED,
      ACOUT(0) => NLW_blk00000918_ACOUT_0_UNCONNECTED,
      CARRYOUT(3) => NLW_blk00000918_CARRYOUT_3_UNCONNECTED,
      CARRYOUT(2) => NLW_blk00000918_CARRYOUT_2_UNCONNECTED,
      CARRYOUT(1) => NLW_blk00000918_CARRYOUT_1_UNCONNECTED,
      CARRYOUT(0) => NLW_blk00000918_CARRYOUT_0_UNCONNECTED
    );
  blk00000919 : DSP48E
    generic map(
      ACASCREG => 2,
      ALUMODEREG => 0,
      AREG => 2,
      AUTORESET_PATTERN_DETECT => FALSE,
      AUTORESET_PATTERN_DETECT_OPTINV => "MATCH",
      A_INPUT => "DIRECT",
      BCASCREG => 2,
      BREG => 2,
      B_INPUT => "DIRECT",
      CARRYINREG => 0,
      CARRYINSELREG => 0,
      CREG => 1,
      MASK => X"000000000000",
      MREG => 1,
      MULTCARRYINREG => 0,
      OPMODEREG => 0,
      PATTERN => X"000000000000",
      PREG => 1,
      SEL_MASK => "MASK",
      SEL_PATTERN => "PATTERN",
      SEL_ROUNDING_MASK => "SEL_MASK",
      SIM_MODE => "SAFE",
      USE_MULT => "MULT_S",
      USE_PATTERN_DETECT => "NO_PATDET",
      USE_SIMD => "ONE48"
    )
    port map (
      CARRYIN => sig000008b6,
      CEA1 => ce,
      CEA2 => ce,
      CEB1 => ce,
      CEB2 => ce,
      CEC => ce,
      CECTRL => sig000008b6,
      CEP => ce,
      CEM => ce,
      CECARRYIN => sig000008b6,
      CEMULTCARRYIN => sig000008b6,
      CLK => clk,
      RSTA => sig000008b6,
      RSTB => sig000008b6,
      RSTC => sig000008b6,
      RSTCTRL => sig000008b6,
      RSTP => sig000008b6,
      RSTM => sig000008b6,
      RSTALLCARRYIN => sig000008b6,
      CEALUMODE => sig000008b6,
      RSTALUMODE => sig000008b6,
      PATTERNBDETECT => NLW_blk00000919_PATTERNBDETECT_UNCONNECTED,
      PATTERNDETECT => NLW_blk00000919_PATTERNDETECT_UNCONNECTED,
      OVERFLOW => NLW_blk00000919_OVERFLOW_UNCONNECTED,
      UNDERFLOW => NLW_blk00000919_UNDERFLOW_UNCONNECTED,
      CARRYCASCIN => sig000008b6,
      CARRYCASCOUT => NLW_blk00000919_CARRYCASCOUT_UNCONNECTED,
      MULTSIGNIN => sig000008b6,
      MULTSIGNOUT => NLW_blk00000919_MULTSIGNOUT_UNCONNECTED,
      A(29) => sig000008b6,
      A(28) => sig000008b6,
      A(27) => sig000008b6,
      A(26) => sig000008b6,
      A(25) => sig000008b6,
      A(24) => sig0000085c,
      A(23) => sig0000085c,
      A(22) => sig0000085c,
      A(21) => sig0000085c,
      A(20) => sig0000085c,
      A(19) => sig0000085c,
      A(18) => sig0000085c,
      A(17) => sig0000085c,
      A(16) => sig0000085c,
      A(15) => sig0000085c,
      A(14) => sig0000085c,
      A(13) => sig0000085c,
      A(12) => sig0000085c,
      A(11) => sig0000085d,
      A(10) => sig0000085e,
      A(9) => sig0000085f,
      A(8) => sig00000860,
      A(7) => sig00000861,
      A(6) => sig00000862,
      A(5) => sig00000863,
      A(4) => sig00000864,
      A(3) => sig00000865,
      A(2) => sig00000866,
      A(1) => sig000008b6,
      A(0) => sig000008b6,
      PCIN(47) => sig000008b6,
      PCIN(46) => sig000008b6,
      PCIN(45) => sig000008b6,
      PCIN(44) => sig000008b6,
      PCIN(43) => sig000008b6,
      PCIN(42) => sig000008b6,
      PCIN(41) => sig000008b6,
      PCIN(40) => sig000008b6,
      PCIN(39) => sig000008b6,
      PCIN(38) => sig000008b6,
      PCIN(37) => sig000008b6,
      PCIN(36) => sig000008b6,
      PCIN(35) => sig000008b6,
      PCIN(34) => sig000008b6,
      PCIN(33) => sig000008b6,
      PCIN(32) => sig000008b6,
      PCIN(31) => sig000008b6,
      PCIN(30) => sig000008b6,
      PCIN(29) => sig000008b6,
      PCIN(28) => sig000008b6,
      PCIN(27) => sig000008b6,
      PCIN(26) => sig000008b6,
      PCIN(25) => sig000008b6,
      PCIN(24) => sig000008b6,
      PCIN(23) => sig000008b6,
      PCIN(22) => sig000008b6,
      PCIN(21) => sig000008b6,
      PCIN(20) => sig000008b6,
      PCIN(19) => sig000008b6,
      PCIN(18) => sig000008b6,
      PCIN(17) => sig000008b6,
      PCIN(16) => sig000008b6,
      PCIN(15) => sig000008b6,
      PCIN(14) => sig000008b6,
      PCIN(13) => sig000008b6,
      PCIN(12) => sig000008b6,
      PCIN(11) => sig000008b6,
      PCIN(10) => sig000008b6,
      PCIN(9) => sig000008b6,
      PCIN(8) => sig000008b6,
      PCIN(7) => sig000008b6,
      PCIN(6) => sig000008b6,
      PCIN(5) => sig000008b6,
      PCIN(4) => sig000008b6,
      PCIN(3) => sig000008b6,
      PCIN(2) => sig000008b6,
      PCIN(1) => sig000008b6,
      PCIN(0) => sig000008b6,
      B(17) => sig0000084e,
      B(16) => sig0000084e,
      B(15) => sig0000084e,
      B(14) => sig0000084e,
      B(13) => sig0000084f,
      B(12) => sig00000850,
      B(11) => sig00000851,
      B(10) => sig00000852,
      B(9) => sig00000853,
      B(8) => sig00000854,
      B(7) => sig00000855,
      B(6) => sig00000856,
      B(5) => sig00000857,
      B(4) => sig00000858,
      B(3) => sig00000859,
      B(2) => sig0000085a,
      B(1) => sig0000085b,
      B(0) => sig00000818,
      C(47) => sig00000832,
      C(46) => sig00000832,
      C(45) => sig00000832,
      C(44) => sig00000832,
      C(43) => sig00000832,
      C(42) => sig00000832,
      C(41) => sig00000832,
      C(40) => sig00000832,
      C(39) => sig00000832,
      C(38) => sig00000832,
      C(37) => sig00000832,
      C(36) => sig00000832,
      C(35) => sig00000832,
      C(34) => sig00000832,
      C(33) => sig00000832,
      C(32) => sig00000832,
      C(31) => sig00000832,
      C(30) => sig00000832,
      C(29) => sig00000832,
      C(28) => sig00000832,
      C(27) => sig00000832,
      C(26) => sig00000833,
      C(25) => sig00000834,
      C(24) => sig00000835,
      C(23) => sig00000836,
      C(22) => sig00000837,
      C(21) => sig00000838,
      C(20) => sig00000839,
      C(19) => sig0000083a,
      C(18) => sig0000083b,
      C(17) => sig0000083c,
      C(16) => sig0000083d,
      C(15) => sig0000083e,
      C(14) => sig0000083f,
      C(13) => sig00000840,
      C(12) => sig00000841,
      C(11) => sig00000842,
      C(10) => sig00000843,
      C(9) => sig00000844,
      C(8) => sig00000845,
      C(7) => sig00000846,
      C(6) => sig00000847,
      C(5) => sig00000848,
      C(4) => sig00000849,
      C(3) => sig0000084a,
      C(2) => sig0000084b,
      C(1) => sig0000084c,
      C(0) => sig0000084d,
      CARRYINSEL(2) => sig000008b6,
      CARRYINSEL(1) => sig000008b6,
      CARRYINSEL(0) => sig000008b6,
      OPMODE(6) => sig000008b6,
      OPMODE(5) => sig000006d1,
      OPMODE(4) => sig000006d1,
      OPMODE(3) => sig000008b6,
      OPMODE(2) => sig000006d1,
      OPMODE(1) => sig000008b6,
      OPMODE(0) => sig000006d1,
      BCIN(17) => sig000008b6,
      BCIN(16) => sig000008b6,
      BCIN(15) => sig000008b6,
      BCIN(14) => sig000008b6,
      BCIN(13) => sig000008b6,
      BCIN(12) => sig000008b6,
      BCIN(11) => sig000008b6,
      BCIN(10) => sig000008b6,
      BCIN(9) => sig000008b6,
      BCIN(8) => sig000008b6,
      BCIN(7) => sig000008b6,
      BCIN(6) => sig000008b6,
      BCIN(5) => sig000008b6,
      BCIN(4) => sig000008b6,
      BCIN(3) => sig000008b6,
      BCIN(2) => sig000008b6,
      BCIN(1) => sig000008b6,
      BCIN(0) => sig000008b6,
      ALUMODE(3) => sig000008b6,
      ALUMODE(2) => sig000008b6,
      ALUMODE(1) => sig000008b6,
      ALUMODE(0) => sig000008b6,
      PCOUT(47) => NLW_blk00000919_PCOUT_47_UNCONNECTED,
      PCOUT(46) => NLW_blk00000919_PCOUT_46_UNCONNECTED,
      PCOUT(45) => NLW_blk00000919_PCOUT_45_UNCONNECTED,
      PCOUT(44) => NLW_blk00000919_PCOUT_44_UNCONNECTED,
      PCOUT(43) => NLW_blk00000919_PCOUT_43_UNCONNECTED,
      PCOUT(42) => NLW_blk00000919_PCOUT_42_UNCONNECTED,
      PCOUT(41) => NLW_blk00000919_PCOUT_41_UNCONNECTED,
      PCOUT(40) => NLW_blk00000919_PCOUT_40_UNCONNECTED,
      PCOUT(39) => NLW_blk00000919_PCOUT_39_UNCONNECTED,
      PCOUT(38) => NLW_blk00000919_PCOUT_38_UNCONNECTED,
      PCOUT(37) => NLW_blk00000919_PCOUT_37_UNCONNECTED,
      PCOUT(36) => NLW_blk00000919_PCOUT_36_UNCONNECTED,
      PCOUT(35) => NLW_blk00000919_PCOUT_35_UNCONNECTED,
      PCOUT(34) => NLW_blk00000919_PCOUT_34_UNCONNECTED,
      PCOUT(33) => NLW_blk00000919_PCOUT_33_UNCONNECTED,
      PCOUT(32) => NLW_blk00000919_PCOUT_32_UNCONNECTED,
      PCOUT(31) => NLW_blk00000919_PCOUT_31_UNCONNECTED,
      PCOUT(30) => NLW_blk00000919_PCOUT_30_UNCONNECTED,
      PCOUT(29) => NLW_blk00000919_PCOUT_29_UNCONNECTED,
      PCOUT(28) => NLW_blk00000919_PCOUT_28_UNCONNECTED,
      PCOUT(27) => NLW_blk00000919_PCOUT_27_UNCONNECTED,
      PCOUT(26) => NLW_blk00000919_PCOUT_26_UNCONNECTED,
      PCOUT(25) => NLW_blk00000919_PCOUT_25_UNCONNECTED,
      PCOUT(24) => NLW_blk00000919_PCOUT_24_UNCONNECTED,
      PCOUT(23) => NLW_blk00000919_PCOUT_23_UNCONNECTED,
      PCOUT(22) => NLW_blk00000919_PCOUT_22_UNCONNECTED,
      PCOUT(21) => NLW_blk00000919_PCOUT_21_UNCONNECTED,
      PCOUT(20) => NLW_blk00000919_PCOUT_20_UNCONNECTED,
      PCOUT(19) => NLW_blk00000919_PCOUT_19_UNCONNECTED,
      PCOUT(18) => NLW_blk00000919_PCOUT_18_UNCONNECTED,
      PCOUT(17) => NLW_blk00000919_PCOUT_17_UNCONNECTED,
      PCOUT(16) => NLW_blk00000919_PCOUT_16_UNCONNECTED,
      PCOUT(15) => NLW_blk00000919_PCOUT_15_UNCONNECTED,
      PCOUT(14) => NLW_blk00000919_PCOUT_14_UNCONNECTED,
      PCOUT(13) => NLW_blk00000919_PCOUT_13_UNCONNECTED,
      PCOUT(12) => NLW_blk00000919_PCOUT_12_UNCONNECTED,
      PCOUT(11) => NLW_blk00000919_PCOUT_11_UNCONNECTED,
      PCOUT(10) => NLW_blk00000919_PCOUT_10_UNCONNECTED,
      PCOUT(9) => NLW_blk00000919_PCOUT_9_UNCONNECTED,
      PCOUT(8) => NLW_blk00000919_PCOUT_8_UNCONNECTED,
      PCOUT(7) => NLW_blk00000919_PCOUT_7_UNCONNECTED,
      PCOUT(6) => NLW_blk00000919_PCOUT_6_UNCONNECTED,
      PCOUT(5) => NLW_blk00000919_PCOUT_5_UNCONNECTED,
      PCOUT(4) => NLW_blk00000919_PCOUT_4_UNCONNECTED,
      PCOUT(3) => NLW_blk00000919_PCOUT_3_UNCONNECTED,
      PCOUT(2) => NLW_blk00000919_PCOUT_2_UNCONNECTED,
      PCOUT(1) => NLW_blk00000919_PCOUT_1_UNCONNECTED,
      PCOUT(0) => NLW_blk00000919_PCOUT_0_UNCONNECTED,
      P(47) => NLW_blk00000919_P_47_UNCONNECTED,
      P(46) => NLW_blk00000919_P_46_UNCONNECTED,
      P(45) => NLW_blk00000919_P_45_UNCONNECTED,
      P(44) => NLW_blk00000919_P_44_UNCONNECTED,
      P(43) => NLW_blk00000919_P_43_UNCONNECTED,
      P(42) => sig000009a5,
      P(41) => sig000009a4,
      P(40) => sig000009a3,
      P(39) => sig000009a2,
      P(38) => sig000009a1,
      P(37) => sig000009a0,
      P(36) => sig0000099f,
      P(35) => sig0000099e,
      P(34) => sig0000099d,
      P(33) => sig0000099c,
      P(32) => sig0000099b,
      P(31) => sig0000099a,
      P(30) => sig00000999,
      P(29) => sig00000998,
      P(28) => sig00000997,
      P(27) => sig00000996,
      P(26) => sig00000995,
      P(25) => sig00000994,
      P(24) => sig00000993,
      P(23) => sig00000992,
      P(22) => sig00000991,
      P(21) => sig00000990,
      P(20) => sig0000098f,
      P(19) => sig0000098e,
      P(18) => sig0000098d,
      P(17) => sig0000098c,
      P(16) => sig0000098b,
      P(15) => sig0000098a,
      P(14) => sig00000989,
      P(13) => sig00000988,
      P(12) => sig00000987,
      P(11) => sig00000986,
      P(10) => sig00000985,
      P(9) => sig00000984,
      P(8) => sig00000983,
      P(7) => sig00000982,
      P(6) => sig00000981,
      P(5) => sig00000980,
      P(4) => sig0000097f,
      P(3) => sig0000097e,
      P(2) => sig0000097d,
      P(1) => sig0000097c,
      P(0) => sig0000097b,
      BCOUT(17) => NLW_blk00000919_BCOUT_17_UNCONNECTED,
      BCOUT(16) => NLW_blk00000919_BCOUT_16_UNCONNECTED,
      BCOUT(15) => NLW_blk00000919_BCOUT_15_UNCONNECTED,
      BCOUT(14) => NLW_blk00000919_BCOUT_14_UNCONNECTED,
      BCOUT(13) => NLW_blk00000919_BCOUT_13_UNCONNECTED,
      BCOUT(12) => NLW_blk00000919_BCOUT_12_UNCONNECTED,
      BCOUT(11) => NLW_blk00000919_BCOUT_11_UNCONNECTED,
      BCOUT(10) => NLW_blk00000919_BCOUT_10_UNCONNECTED,
      BCOUT(9) => NLW_blk00000919_BCOUT_9_UNCONNECTED,
      BCOUT(8) => NLW_blk00000919_BCOUT_8_UNCONNECTED,
      BCOUT(7) => NLW_blk00000919_BCOUT_7_UNCONNECTED,
      BCOUT(6) => NLW_blk00000919_BCOUT_6_UNCONNECTED,
      BCOUT(5) => NLW_blk00000919_BCOUT_5_UNCONNECTED,
      BCOUT(4) => NLW_blk00000919_BCOUT_4_UNCONNECTED,
      BCOUT(3) => NLW_blk00000919_BCOUT_3_UNCONNECTED,
      BCOUT(2) => NLW_blk00000919_BCOUT_2_UNCONNECTED,
      BCOUT(1) => NLW_blk00000919_BCOUT_1_UNCONNECTED,
      BCOUT(0) => NLW_blk00000919_BCOUT_0_UNCONNECTED,
      ACIN(29) => sig000008b6,
      ACIN(28) => sig000008b6,
      ACIN(27) => sig000008b6,
      ACIN(26) => sig000008b6,
      ACIN(25) => sig000008b6,
      ACIN(24) => sig000008b6,
      ACIN(23) => sig000008b6,
      ACIN(22) => sig000008b6,
      ACIN(21) => sig000008b6,
      ACIN(20) => sig000008b6,
      ACIN(19) => sig000008b6,
      ACIN(18) => sig000008b6,
      ACIN(17) => sig000008b6,
      ACIN(16) => sig000008b6,
      ACIN(15) => sig000008b6,
      ACIN(14) => sig000008b6,
      ACIN(13) => sig000008b6,
      ACIN(12) => sig000008b6,
      ACIN(11) => sig000008b6,
      ACIN(10) => sig000008b6,
      ACIN(9) => sig000008b6,
      ACIN(8) => sig000008b6,
      ACIN(7) => sig000008b6,
      ACIN(6) => sig000008b6,
      ACIN(5) => sig000008b6,
      ACIN(4) => sig000008b6,
      ACIN(3) => sig000008b6,
      ACIN(2) => sig000008b6,
      ACIN(1) => sig000008b6,
      ACIN(0) => sig000008b6,
      ACOUT(29) => NLW_blk00000919_ACOUT_29_UNCONNECTED,
      ACOUT(28) => NLW_blk00000919_ACOUT_28_UNCONNECTED,
      ACOUT(27) => NLW_blk00000919_ACOUT_27_UNCONNECTED,
      ACOUT(26) => NLW_blk00000919_ACOUT_26_UNCONNECTED,
      ACOUT(25) => NLW_blk00000919_ACOUT_25_UNCONNECTED,
      ACOUT(24) => NLW_blk00000919_ACOUT_24_UNCONNECTED,
      ACOUT(23) => NLW_blk00000919_ACOUT_23_UNCONNECTED,
      ACOUT(22) => NLW_blk00000919_ACOUT_22_UNCONNECTED,
      ACOUT(21) => NLW_blk00000919_ACOUT_21_UNCONNECTED,
      ACOUT(20) => NLW_blk00000919_ACOUT_20_UNCONNECTED,
      ACOUT(19) => NLW_blk00000919_ACOUT_19_UNCONNECTED,
      ACOUT(18) => NLW_blk00000919_ACOUT_18_UNCONNECTED,
      ACOUT(17) => NLW_blk00000919_ACOUT_17_UNCONNECTED,
      ACOUT(16) => NLW_blk00000919_ACOUT_16_UNCONNECTED,
      ACOUT(15) => NLW_blk00000919_ACOUT_15_UNCONNECTED,
      ACOUT(14) => NLW_blk00000919_ACOUT_14_UNCONNECTED,
      ACOUT(13) => NLW_blk00000919_ACOUT_13_UNCONNECTED,
      ACOUT(12) => NLW_blk00000919_ACOUT_12_UNCONNECTED,
      ACOUT(11) => NLW_blk00000919_ACOUT_11_UNCONNECTED,
      ACOUT(10) => NLW_blk00000919_ACOUT_10_UNCONNECTED,
      ACOUT(9) => NLW_blk00000919_ACOUT_9_UNCONNECTED,
      ACOUT(8) => NLW_blk00000919_ACOUT_8_UNCONNECTED,
      ACOUT(7) => NLW_blk00000919_ACOUT_7_UNCONNECTED,
      ACOUT(6) => NLW_blk00000919_ACOUT_6_UNCONNECTED,
      ACOUT(5) => NLW_blk00000919_ACOUT_5_UNCONNECTED,
      ACOUT(4) => NLW_blk00000919_ACOUT_4_UNCONNECTED,
      ACOUT(3) => NLW_blk00000919_ACOUT_3_UNCONNECTED,
      ACOUT(2) => NLW_blk00000919_ACOUT_2_UNCONNECTED,
      ACOUT(1) => NLW_blk00000919_ACOUT_1_UNCONNECTED,
      ACOUT(0) => NLW_blk00000919_ACOUT_0_UNCONNECTED,
      CARRYOUT(3) => NLW_blk00000919_CARRYOUT_3_UNCONNECTED,
      CARRYOUT(2) => NLW_blk00000919_CARRYOUT_2_UNCONNECTED,
      CARRYOUT(1) => NLW_blk00000919_CARRYOUT_1_UNCONNECTED,
      CARRYOUT(0) => NLW_blk00000919_CARRYOUT_0_UNCONNECTED
    );
  blk00000920 : FDR
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      D => sig000009f6,
      R => sig000008b6,
      Q => sig000000ca
    );
  blk00000921 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => sig000009f8,
      D => sig0000010d,
      Q => sig00000a5b
    );
  blk00000922 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => sig000009f8,
      D => sig0000010e,
      Q => sig00000a5c
    );
  blk00000923 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => sig000009f8,
      D => sig0000010f,
      Q => sig00000a5d
    );
  blk00000924 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => sig000009f8,
      D => sig00000110,
      Q => sig00000a5e
    );
  blk00000925 : FD
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      D => sig000009f7,
      Q => sig00000a60
    );
  blk00000926 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => sig000009f8,
      D => sig00000a60,
      Q => sig000009f9
    );
  blk00000927 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => sig000009f8,
      D => sig0000010c,
      Q => sig00000a66
    );
  blk00000928 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => sig000009f8,
      D => sig0000010b,
      Q => sig00000a65
    );
  blk00000929 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => sig000009f8,
      D => sig0000010a,
      Q => sig00000a64
    );
  blk0000092a : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => sig000009f8,
      D => sig00000109,
      Q => sig00000a63
    );
  blk0000092b : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => sig000009f8,
      D => sig00000108,
      Q => sig00000a62
    );
  blk0000092c : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => sig000009f8,
      D => sig00000107,
      Q => sig00000a61
    );
  blk00000944 : LUT6
    generic map(
      INIT => X"9009000000009009"
    )
    port map (
      I0 => sig00000a8a,
      I1 => sig000008b6,
      I2 => sig00000aa3,
      I3 => sig000008b6,
      I4 => sig00000aa4,
      I5 => sig000008b6,
      O => sig00000a8b
    );
  blk00000945 : LUT6
    generic map(
      INIT => X"9009000000009009"
    )
    port map (
      I0 => sig00000a87,
      I1 => sig000008b6,
      I2 => sig00000a88,
      I3 => sig000006d1,
      I4 => sig00000a89,
      I5 => sig000008b6,
      O => sig00000a8c
    );
  blk00000946 : MUXCY
    port map (
      CI => sig00000a8d,
      DI => sig000008b6,
      S => sig00000a8b,
      O => sig00000a9e
    );
  blk00000947 : MUXCY
    port map (
      CI => sig000006d1,
      DI => sig000008b6,
      S => sig00000a8c,
      O => sig00000a8d
    );
  blk00000948 : LUT6
    generic map(
      INIT => X"9009000000009009"
    )
    port map (
      I0 => sig00000a8a,
      I1 => sig000006d1,
      I2 => sig00000aa3,
      I3 => sig000006d1,
      I4 => sig00000aa4,
      I5 => sig000006d1,
      O => sig00000a8e
    );
  blk00000949 : LUT6
    generic map(
      INIT => X"9009000000009009"
    )
    port map (
      I0 => sig00000a87,
      I1 => sig000006d1,
      I2 => sig00000a88,
      I3 => sig000008b6,
      I4 => sig00000a89,
      I5 => sig000006d1,
      O => sig00000a8f
    );
  blk0000094a : MUXCY
    port map (
      CI => sig00000a91,
      DI => sig000008b6,
      S => sig00000a8e,
      O => sig00000a90
    );
  blk0000094b : MUXCY
    port map (
      CI => sig000006d1,
      DI => sig000008b6,
      S => sig00000a8f,
      O => sig00000a91
    );
  blk0000094c : XORCY
    port map (
      CI => sig00000a90,
      LI => sig000008b6,
      O => sig00000a92
    );
  blk0000094d : MUXCY
    port map (
      CI => sig000006d1,
      DI => sig000008b6,
      S => sig00000a9a,
      O => sig00000a9b
    );
  blk0000094e : XORCY
    port map (
      CI => sig00000a9d,
      LI => sig000008b6,
      O => sig00000a9c
    );
  blk0000094f : MUXCY
    port map (
      CI => sig00000a9e,
      DI => sig000008b6,
      S => sig00000aa0,
      O => sig00000a9d
    );
  blk00000950 : LUT3
    generic map(
      INIT => X"AE"
    )
    port map (
      I0 => sig000000ee,
      I1 => sig00000aa1,
      I2 => sig00000aa2,
      O => sig00000a9f
    );
  blk00000951 : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => sig00000aa0,
      D => sig00000a93,
      R => sig000008b6,
      Q => sig00000aa2
    );
  blk00000952 : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => sig00000aa0,
      D => sig00000a92,
      R => sig000008b6,
      Q => sig00000a93
    );
  blk00000953 : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => sig00000a9c,
      R => sig000008b6,
      Q => sig00000a86
    );
  blk00000954 : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => sig00000a9f,
      R => sig000008b6,
      Q => sig00000aa1
    );
  blk0000096c : LUT6
    generic map(
      INIT => X"9009000000009009"
    )
    port map (
      I0 => sig00000a85,
      I1 => sig000008b6,
      I2 => sig00000abd,
      I3 => sig000008b6,
      I4 => sig00000abe,
      I5 => sig000008b6,
      O => sig00000aa5
    );
  blk0000096d : LUT6
    generic map(
      INIT => X"9009000000009009"
    )
    port map (
      I0 => sig00000a82,
      I1 => sig000008b6,
      I2 => sig00000a83,
      I3 => sig000008b6,
      I4 => sig00000a84,
      I5 => sig000008b6,
      O => sig00000aa6
    );
  blk0000096e : MUXCY
    port map (
      CI => sig00000aa7,
      DI => sig000008b6,
      S => sig00000aa5,
      O => sig00000ab8
    );
  blk0000096f : MUXCY
    port map (
      CI => sig000006d1,
      DI => sig000008b6,
      S => sig00000aa6,
      O => sig00000aa7
    );
  blk00000970 : LUT6
    generic map(
      INIT => X"9009000000009009"
    )
    port map (
      I0 => sig00000a85,
      I1 => sig000006d1,
      I2 => sig00000abd,
      I3 => sig000006d1,
      I4 => sig00000abe,
      I5 => sig000006d1,
      O => sig00000aa8
    );
  blk00000971 : LUT6
    generic map(
      INIT => X"9009000000009009"
    )
    port map (
      I0 => sig00000a82,
      I1 => sig000006d1,
      I2 => sig00000a83,
      I3 => sig000008b6,
      I4 => sig00000a84,
      I5 => sig000006d1,
      O => sig00000aa9
    );
  blk00000972 : MUXCY
    port map (
      CI => sig00000aab,
      DI => sig000008b6,
      S => sig00000aa8,
      O => sig00000aaa
    );
  blk00000973 : MUXCY
    port map (
      CI => sig000006d1,
      DI => sig000008b6,
      S => sig00000aa9,
      O => sig00000aab
    );
  blk00000974 : XORCY
    port map (
      CI => sig00000aaa,
      LI => sig000008b6,
      O => sig00000aac
    );
  blk00000975 : MUXCY
    port map (
      CI => sig000006d1,
      DI => sig000008b6,
      S => sig00000ab4,
      O => sig00000ab5
    );
  blk00000976 : XORCY
    port map (
      CI => sig00000ab7,
      LI => sig000008b6,
      O => sig00000ab6
    );
  blk00000977 : MUXCY
    port map (
      CI => sig00000ab8,
      DI => sig000008b6,
      S => sig00000aba,
      O => sig00000ab7
    );
  blk00000978 : LUT3
    generic map(
      INIT => X"AE"
    )
    port map (
      I0 => sig00000a86,
      I1 => sig00000abb,
      I2 => sig00000abc,
      O => sig00000ab9
    );
  blk00000979 : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => sig00000aba,
      D => sig00000aad,
      R => sig000008b6,
      Q => sig00000abc
    );
  blk0000097a : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => sig00000aba,
      D => sig00000aac,
      R => sig000008b6,
      Q => sig00000aad
    );
  blk0000097b : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => sig00000ab6,
      R => sig000008b6,
      Q => sig00000a81
    );
  blk0000097c : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => sig00000ab9,
      R => sig000008b6,
      Q => sig00000abb
    );
  blk0000097d : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => sig00000acb,
      R => sig000008b6,
      Q => sig00000af1
    );
  blk0000097e : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => sig00000aca,
      R => sig000008b6,
      Q => sig00000af2
    );
  blk0000097f : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => sig00000ac9,
      R => sig000008b6,
      Q => sig00000af3
    );
  blk00000980 : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => sig00000ac8,
      R => sig000008b6,
      Q => sig00000af4
    );
  blk00000981 : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => sig00000ac7,
      R => sig000008b6,
      Q => sig00000af5
    );
  blk00000982 : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => sig00000ac6,
      R => sig000008b6,
      Q => sig00000af6
    );
  blk00000983 : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => sig00000ac5,
      R => sig000008b6,
      Q => sig00000af7
    );
  blk00000984 : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => sig00000ac4,
      R => sig000008b6,
      Q => sig00000af8
    );
  blk00000985 : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => sig00000ac3,
      R => sig000008b6,
      Q => sig00000af9
    );
  blk00000986 : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => sig00000ac2,
      R => sig000008b6,
      Q => sig00000afa
    );
  blk00000987 : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => sig00000ac1,
      R => sig000008b6,
      Q => sig00000afb
    );
  blk00000988 : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => sig00000ac0,
      R => sig000008b6,
      Q => sig00000afc
    );
  blk00000989 : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => sig00000abf,
      R => sig000008b6,
      Q => sig00000afd
    );
  blk0000098a : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => sig00000ad8,
      R => sig000008b6,
      Q => sig00000a67
    );
  blk0000098b : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => sig00000ad7,
      R => sig000008b6,
      Q => sig00000a68
    );
  blk0000098c : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => sig00000ad6,
      R => sig000008b6,
      Q => sig00000a69
    );
  blk0000098d : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => sig00000ad5,
      R => sig000008b6,
      Q => sig00000a6a
    );
  blk0000098e : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => sig00000ad4,
      R => sig000008b6,
      Q => sig00000a6b
    );
  blk0000098f : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => sig00000ad3,
      R => sig000008b6,
      Q => sig00000a6c
    );
  blk00000990 : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => sig00000ad2,
      R => sig000008b6,
      Q => sig00000a6d
    );
  blk00000991 : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => sig00000ad1,
      R => sig000008b6,
      Q => sig00000a6e
    );
  blk00000992 : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => sig00000ad0,
      R => sig000008b6,
      Q => sig00000a6f
    );
  blk00000993 : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => sig00000acf,
      R => sig000008b6,
      Q => sig00000a70
    );
  blk00000994 : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => sig00000ace,
      R => sig000008b6,
      Q => sig00000a71
    );
  blk00000995 : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => sig00000acd,
      R => sig000008b6,
      Q => sig00000a72
    );
  blk00000996 : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => sig00000acc,
      R => sig000008b6,
      Q => sig00000a73
    );
  blk00000997 : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => sig00000ae4,
      R => sig000008b6,
      Q => sig00000b4c
    );
  blk00000998 : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => sig00000ae3,
      R => sig000008b6,
      Q => sig00000b4d
    );
  blk00000999 : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => sig00000ae2,
      R => sig000008b6,
      Q => sig00000b4e
    );
  blk0000099a : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => sig00000ae1,
      R => sig000008b6,
      Q => sig00000b4f
    );
  blk0000099b : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => sig00000ae0,
      R => sig000008b6,
      Q => sig00000b50
    );
  blk0000099c : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => sig00000adf,
      R => sig000008b6,
      Q => sig00000b51
    );
  blk0000099d : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => sig00000ade,
      R => sig000008b6,
      Q => sig00000b52
    );
  blk0000099e : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => sig00000add,
      R => sig000008b6,
      Q => sig00000b53
    );
  blk0000099f : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => sig00000adc,
      R => sig000008b6,
      Q => sig00000b54
    );
  blk000009a0 : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => sig00000adb,
      R => sig000008b6,
      Q => sig00000b55
    );
  blk000009a1 : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => sig00000ada,
      R => sig000008b6,
      Q => sig00000b56
    );
  blk000009a2 : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => sig00000ad9,
      R => sig000008b6,
      Q => sig00000b57
    );
  blk000009a3 : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => sig00000af0,
      R => sig000008b6,
      Q => sig00000b40
    );
  blk000009a4 : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => sig00000aef,
      R => sig000008b6,
      Q => sig00000b41
    );
  blk000009a5 : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => sig00000aee,
      R => sig000008b6,
      Q => sig00000b42
    );
  blk000009a6 : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => sig00000aed,
      R => sig000008b6,
      Q => sig00000b43
    );
  blk000009a7 : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => sig00000aec,
      R => sig000008b6,
      Q => sig00000b44
    );
  blk000009a8 : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => sig00000aeb,
      R => sig000008b6,
      Q => sig00000b45
    );
  blk000009a9 : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => sig00000aea,
      R => sig000008b6,
      Q => sig00000b46
    );
  blk000009aa : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => sig00000ae9,
      R => sig000008b6,
      Q => sig00000b47
    );
  blk000009ab : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => sig00000ae8,
      R => sig000008b6,
      Q => sig00000b48
    );
  blk000009ac : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => sig00000ae7,
      R => sig000008b6,
      Q => sig00000b49
    );
  blk000009ad : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => sig00000ae6,
      R => sig000008b6,
      Q => sig00000b4a
    );
  blk000009ae : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => sig00000ae5,
      R => sig000008b6,
      Q => sig00000b4b
    );
  blk000009af : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => sig00000b33,
      Q => sig00000b32
    );
  blk000009b0 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => sig00000111,
      Q => sig00000b33
    );
  blk00000b59 : MUXCY
    port map (
      CI => sig00000bb9,
      DI => sig000008b6,
      S => sig00000b90,
      O => sig00000b9e
    );
  blk00000b5a : XORCY
    port map (
      CI => sig00000bb9,
      LI => sig00000b90,
      O => sig00000b9f
    );
  blk00000b5b : MUXCY
    port map (
      CI => sig00000b9e,
      DI => sig000008b6,
      S => sig00000b91,
      O => sig00000ba0
    );
  blk00000b5c : XORCY
    port map (
      CI => sig00000b9e,
      LI => sig00000b91,
      O => sig00000ba1
    );
  blk00000b5d : MUXCY
    port map (
      CI => sig00000ba0,
      DI => sig000008b6,
      S => sig00000b92,
      O => sig00000ba2
    );
  blk00000b5e : XORCY
    port map (
      CI => sig00000ba0,
      LI => sig00000b92,
      O => sig00000ba3
    );
  blk00000b5f : MUXCY
    port map (
      CI => sig00000ba2,
      DI => sig000008b6,
      S => sig00000b93,
      O => sig00000ba4
    );
  blk00000b60 : XORCY
    port map (
      CI => sig00000ba2,
      LI => sig00000b93,
      O => sig00000ba5
    );
  blk00000b61 : MUXCY
    port map (
      CI => sig00000ba4,
      DI => sig000008b6,
      S => sig00000b94,
      O => sig00000ba6
    );
  blk00000b62 : XORCY
    port map (
      CI => sig00000ba4,
      LI => sig00000b94,
      O => sig00000ba7
    );
  blk00000b63 : MUXCY
    port map (
      CI => sig00000ba6,
      DI => sig000008b6,
      S => sig00000b95,
      O => sig00000ba8
    );
  blk00000b64 : XORCY
    port map (
      CI => sig00000ba6,
      LI => sig00000b95,
      O => sig00000ba9
    );
  blk00000b65 : MUXCY
    port map (
      CI => sig00000ba8,
      DI => sig000008b6,
      S => sig00000b96,
      O => sig00000baa
    );
  blk00000b66 : XORCY
    port map (
      CI => sig00000ba8,
      LI => sig00000b96,
      O => sig00000bab
    );
  blk00000b67 : MUXCY
    port map (
      CI => sig00000baa,
      DI => sig000008b6,
      S => sig00000b97,
      O => sig00000bac
    );
  blk00000b68 : XORCY
    port map (
      CI => sig00000baa,
      LI => sig00000b97,
      O => sig00000bad
    );
  blk00000b69 : MUXCY
    port map (
      CI => sig00000bac,
      DI => sig000008b6,
      S => sig00000b98,
      O => sig00000bae
    );
  blk00000b6a : XORCY
    port map (
      CI => sig00000bac,
      LI => sig00000b98,
      O => sig00000baf
    );
  blk00000b6b : MUXCY
    port map (
      CI => sig00000bae,
      DI => sig000008b6,
      S => sig00000b99,
      O => sig00000bb0
    );
  blk00000b6c : XORCY
    port map (
      CI => sig00000bae,
      LI => sig00000b99,
      O => sig00000bb1
    );
  blk00000b6d : MUXCY
    port map (
      CI => sig00000bb0,
      DI => sig000008b6,
      S => sig00000b9a,
      O => sig00000bb2
    );
  blk00000b6e : XORCY
    port map (
      CI => sig00000bb0,
      LI => sig00000b9a,
      O => sig00000bb3
    );
  blk00000b6f : MUXCY
    port map (
      CI => sig00000bb2,
      DI => sig000008b6,
      S => sig00000b9b,
      O => sig00000bb4
    );
  blk00000b70 : XORCY
    port map (
      CI => sig00000bb2,
      LI => sig00000b9b,
      O => sig00000bb5
    );
  blk00000b71 : MUXCY
    port map (
      CI => sig00000bb4,
      DI => sig000008b6,
      S => sig00000ef3,
      O => sig00000bb6
    );
  blk00000b72 : XORCY
    port map (
      CI => sig00000bb4,
      LI => sig00000ef3,
      O => sig00000bb7
    );
  blk00000b73 : MUXCY
    port map (
      CI => sig00000bb6,
      DI => sig000008b6,
      S => sig00000b9c,
      O => NLW_blk00000b73_O_UNCONNECTED
    );
  blk00000b74 : XORCY
    port map (
      CI => sig00000bb6,
      LI => sig00000b9c,
      O => sig00000bb8
    );
  blk00000b75 : MUXCY
    port map (
      CI => sig000006d1,
      DI => sig000008b6,
      S => sig00000b9d,
      O => sig00000bb9
    );
  blk00000b76 : MUXCY
    port map (
      CI => sig00000be3,
      DI => sig000008b6,
      S => sig00000bba,
      O => sig00000bc8
    );
  blk00000b77 : XORCY
    port map (
      CI => sig00000be3,
      LI => sig00000bba,
      O => sig00000bc9
    );
  blk00000b78 : MUXCY
    port map (
      CI => sig00000bc8,
      DI => sig000008b6,
      S => sig00000bbb,
      O => sig00000bca
    );
  blk00000b79 : XORCY
    port map (
      CI => sig00000bc8,
      LI => sig00000bbb,
      O => sig00000bcb
    );
  blk00000b7a : MUXCY
    port map (
      CI => sig00000bca,
      DI => sig000008b6,
      S => sig00000bbc,
      O => sig00000bcc
    );
  blk00000b7b : XORCY
    port map (
      CI => sig00000bca,
      LI => sig00000bbc,
      O => sig00000bcd
    );
  blk00000b7c : MUXCY
    port map (
      CI => sig00000bcc,
      DI => sig000008b6,
      S => sig00000bbd,
      O => sig00000bce
    );
  blk00000b7d : XORCY
    port map (
      CI => sig00000bcc,
      LI => sig00000bbd,
      O => sig00000bcf
    );
  blk00000b7e : MUXCY
    port map (
      CI => sig00000bce,
      DI => sig000008b6,
      S => sig00000bbe,
      O => sig00000bd0
    );
  blk00000b7f : XORCY
    port map (
      CI => sig00000bce,
      LI => sig00000bbe,
      O => sig00000bd1
    );
  blk00000b80 : MUXCY
    port map (
      CI => sig00000bd0,
      DI => sig000008b6,
      S => sig00000bbf,
      O => sig00000bd2
    );
  blk00000b81 : XORCY
    port map (
      CI => sig00000bd0,
      LI => sig00000bbf,
      O => sig00000bd3
    );
  blk00000b82 : MUXCY
    port map (
      CI => sig00000bd2,
      DI => sig000008b6,
      S => sig00000bc0,
      O => sig00000bd4
    );
  blk00000b83 : XORCY
    port map (
      CI => sig00000bd2,
      LI => sig00000bc0,
      O => sig00000bd5
    );
  blk00000b84 : MUXCY
    port map (
      CI => sig00000bd4,
      DI => sig000008b6,
      S => sig00000bc1,
      O => sig00000bd6
    );
  blk00000b85 : XORCY
    port map (
      CI => sig00000bd4,
      LI => sig00000bc1,
      O => sig00000bd7
    );
  blk00000b86 : MUXCY
    port map (
      CI => sig00000bd6,
      DI => sig000008b6,
      S => sig00000bc2,
      O => sig00000bd8
    );
  blk00000b87 : XORCY
    port map (
      CI => sig00000bd6,
      LI => sig00000bc2,
      O => sig00000bd9
    );
  blk00000b88 : MUXCY
    port map (
      CI => sig00000bd8,
      DI => sig000008b6,
      S => sig00000bc3,
      O => sig00000bda
    );
  blk00000b89 : XORCY
    port map (
      CI => sig00000bd8,
      LI => sig00000bc3,
      O => sig00000bdb
    );
  blk00000b8a : MUXCY
    port map (
      CI => sig00000bda,
      DI => sig000008b6,
      S => sig00000bc4,
      O => sig00000bdc
    );
  blk00000b8b : XORCY
    port map (
      CI => sig00000bda,
      LI => sig00000bc4,
      O => sig00000bdd
    );
  blk00000b8c : MUXCY
    port map (
      CI => sig00000bdc,
      DI => sig000008b6,
      S => sig00000bc5,
      O => sig00000bde
    );
  blk00000b8d : XORCY
    port map (
      CI => sig00000bdc,
      LI => sig00000bc5,
      O => sig00000bdf
    );
  blk00000b8e : MUXCY
    port map (
      CI => sig00000bde,
      DI => sig000008b6,
      S => sig00000ef4,
      O => sig00000be0
    );
  blk00000b8f : XORCY
    port map (
      CI => sig00000bde,
      LI => sig00000ef4,
      O => sig00000be1
    );
  blk00000b90 : MUXCY
    port map (
      CI => sig00000be0,
      DI => sig000008b6,
      S => sig00000bc6,
      O => NLW_blk00000b90_O_UNCONNECTED
    );
  blk00000b91 : XORCY
    port map (
      CI => sig00000be0,
      LI => sig00000bc6,
      O => sig00000be2
    );
  blk00000b92 : MUXCY
    port map (
      CI => sig000006d1,
      DI => sig000008b6,
      S => sig00000bc7,
      O => sig00000be3
    );
  blk00000b93 : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => sig00000b65,
      R => sig000008b6,
      Q => sig00000c47
    );
  blk00000b94 : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => sig00000b64,
      R => sig000008b6,
      Q => sig00000c48
    );
  blk00000b95 : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => sig00000b63,
      R => sig000008b6,
      Q => sig00000c49
    );
  blk00000b96 : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => sig00000b62,
      R => sig000008b6,
      Q => sig00000c4a
    );
  blk00000b97 : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => sig00000b61,
      R => sig000008b6,
      Q => sig00000c4b
    );
  blk00000b98 : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => sig00000b60,
      R => sig000008b6,
      Q => sig00000c4c
    );
  blk00000b99 : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => sig00000b5f,
      R => sig000008b6,
      Q => sig00000c4d
    );
  blk00000b9a : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => sig00000b5e,
      R => sig000008b6,
      Q => sig00000c4e
    );
  blk00000b9b : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => sig00000b5d,
      R => sig000008b6,
      Q => sig00000c4f
    );
  blk00000b9c : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => sig00000b5c,
      R => sig000008b6,
      Q => sig00000c50
    );
  blk00000b9d : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => sig00000b5b,
      R => sig000008b6,
      Q => sig00000c51
    );
  blk00000b9e : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => sig00000b5a,
      R => sig000008b6,
      Q => sig00000c52
    );
  blk00000b9f : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => sig00000b59,
      R => sig000008b6,
      Q => sig00000c53
    );
  blk00000ba0 : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => sig00000b58,
      R => sig000008b6,
      Q => sig00000c54
    );
  blk00000ba1 : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => sig00000b73,
      R => sig000008b6,
      Q => sig00000c39
    );
  blk00000ba2 : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => sig00000b72,
      R => sig000008b6,
      Q => sig00000c3a
    );
  blk00000ba3 : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => sig00000b71,
      R => sig000008b6,
      Q => sig00000c3b
    );
  blk00000ba4 : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => sig00000b70,
      R => sig000008b6,
      Q => sig00000c3c
    );
  blk00000ba5 : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => sig00000b6f,
      R => sig000008b6,
      Q => sig00000c3d
    );
  blk00000ba6 : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => sig00000b6e,
      R => sig000008b6,
      Q => sig00000c3e
    );
  blk00000ba7 : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => sig00000b6d,
      R => sig000008b6,
      Q => sig00000c3f
    );
  blk00000ba8 : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => sig00000b6c,
      R => sig000008b6,
      Q => sig00000c40
    );
  blk00000ba9 : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => sig00000b6b,
      R => sig000008b6,
      Q => sig00000c41
    );
  blk00000baa : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => sig00000b6a,
      R => sig000008b6,
      Q => sig00000c42
    );
  blk00000bab : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => sig00000b69,
      R => sig000008b6,
      Q => sig00000c43
    );
  blk00000bac : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => sig00000b68,
      R => sig000008b6,
      Q => sig00000c44
    );
  blk00000bad : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => sig00000b67,
      R => sig000008b6,
      Q => sig00000c45
    );
  blk00000bae : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => sig00000b66,
      R => sig000008b6,
      Q => sig00000c46
    );
  blk00000baf : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => sig00000b81,
      R => sig000008b6,
      Q => sig00000c01
    );
  blk00000bb0 : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => sig00000b80,
      R => sig000008b6,
      Q => sig00000c02
    );
  blk00000bb1 : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => sig00000b7f,
      R => sig000008b6,
      Q => sig00000c03
    );
  blk00000bb2 : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => sig00000b7e,
      R => sig000008b6,
      Q => sig00000c04
    );
  blk00000bb3 : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => sig00000b7d,
      R => sig000008b6,
      Q => sig00000c05
    );
  blk00000bb4 : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => sig00000b7c,
      R => sig000008b6,
      Q => sig00000c06
    );
  blk00000bb5 : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => sig00000b7b,
      R => sig000008b6,
      Q => sig00000c07
    );
  blk00000bb6 : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => sig00000b7a,
      R => sig000008b6,
      Q => sig00000c08
    );
  blk00000bb7 : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => sig00000b79,
      R => sig000008b6,
      Q => sig00000c09
    );
  blk00000bb8 : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => sig00000b78,
      R => sig000008b6,
      Q => sig00000c0a
    );
  blk00000bb9 : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => sig00000b77,
      R => sig000008b6,
      Q => sig00000c0b
    );
  blk00000bba : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => sig00000b76,
      R => sig000008b6,
      Q => sig00000c0c
    );
  blk00000bbb : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => sig00000b75,
      R => sig000008b6,
      Q => sig00000c0d
    );
  blk00000bbc : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => sig00000b74,
      R => sig000008b6,
      Q => sig00000c0e
    );
  blk00000bbd : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => sig00000b8f,
      R => sig000008b6,
      Q => sig00000a3b
    );
  blk00000bbe : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => sig00000b8e,
      R => sig000008b6,
      Q => sig00000a3c
    );
  blk00000bbf : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => sig00000b8d,
      R => sig000008b6,
      Q => sig00000a3d
    );
  blk00000bc0 : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => sig00000b8c,
      R => sig000008b6,
      Q => sig00000a3e
    );
  blk00000bc1 : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => sig00000b8b,
      R => sig000008b6,
      Q => sig00000a3f
    );
  blk00000bc2 : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => sig00000b8a,
      R => sig000008b6,
      Q => sig00000a40
    );
  blk00000bc3 : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => sig00000b89,
      R => sig000008b6,
      Q => sig00000a41
    );
  blk00000bc4 : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => sig00000b88,
      R => sig000008b6,
      Q => sig00000a42
    );
  blk00000bc5 : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => sig00000b87,
      R => sig000008b6,
      Q => sig00000a43
    );
  blk00000bc6 : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => sig00000b86,
      R => sig000008b6,
      Q => sig00000a44
    );
  blk00000bc7 : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => sig00000b85,
      R => sig000008b6,
      Q => sig00000a45
    );
  blk00000bc8 : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => sig00000b84,
      R => sig000008b6,
      Q => sig00000a46
    );
  blk00000bc9 : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => sig00000b83,
      R => sig000008b6,
      Q => sig00000a47
    );
  blk00000bca : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => sig00000b82,
      R => sig000008b6,
      Q => sig00000a48
    );
  blk00000bcb : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => sig00000b9f,
      Q => sig00000c71
    );
  blk00000bcc : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => sig00000ba1,
      Q => sig00000c72
    );
  blk00000bcd : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => sig00000ba3,
      Q => sig00000c73
    );
  blk00000bce : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => sig00000ba5,
      Q => sig00000c74
    );
  blk00000bcf : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => sig00000ba7,
      Q => sig00000c75
    );
  blk00000bd0 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => sig00000ba9,
      Q => sig00000c76
    );
  blk00000bd1 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => sig00000bab,
      Q => sig00000c77
    );
  blk00000bd2 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => sig00000bad,
      Q => sig00000c78
    );
  blk00000bd3 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => sig00000baf,
      Q => sig00000c79
    );
  blk00000bd4 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => sig00000bb1,
      Q => sig00000c7a
    );
  blk00000bd5 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => sig00000bb3,
      Q => sig00000c7b
    );
  blk00000bd6 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => sig00000bb5,
      Q => sig00000c7c
    );
  blk00000bd7 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => sig00000bb7,
      Q => sig00000c7d
    );
  blk00000bd8 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => sig00000bb8,
      Q => sig00000c7e
    );
  blk00000bd9 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => sig00000bc9,
      Q => sig00000c7f
    );
  blk00000bda : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => sig00000bcb,
      Q => sig00000c80
    );
  blk00000bdb : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => sig00000bcd,
      Q => sig00000c81
    );
  blk00000bdc : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => sig00000bcf,
      Q => sig00000c82
    );
  blk00000bdd : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => sig00000bd1,
      Q => sig00000c83
    );
  blk00000bde : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => sig00000bd3,
      Q => sig00000c84
    );
  blk00000bdf : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => sig00000bd5,
      Q => sig00000c85
    );
  blk00000be0 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => sig00000bd7,
      Q => sig00000c86
    );
  blk00000be1 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => sig00000bd9,
      Q => sig00000c87
    );
  blk00000be2 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => sig00000bdb,
      Q => sig00000c88
    );
  blk00000be3 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => sig00000bdd,
      Q => sig00000c89
    );
  blk00000be4 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => sig00000bdf,
      Q => sig00000c8a
    );
  blk00000be5 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => sig00000be1,
      Q => sig00000c8b
    );
  blk00000be6 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => sig00000be2,
      Q => sig00000c8c
    );
  blk00000be7 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => sig00000a5f,
      Q => sig00000c92
    );
  blk00000be8 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => sig00000be4,
      Q => sig00000c8d
    );
  blk00000be9 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => sig00000a57,
      Q => sig00000c91
    );
  blk00000bea : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => sig00000c8c,
      Q => sig00000bf2
    );
  blk00000beb : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => sig00000c8b,
      Q => sig00000bf1
    );
  blk00000bec : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => sig00000c8a,
      Q => sig00000bf0
    );
  blk00000bed : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => sig00000c89,
      Q => sig00000bef
    );
  blk00000bee : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => sig00000c88,
      Q => sig00000bee
    );
  blk00000bef : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => sig00000c87,
      Q => sig00000bed
    );
  blk00000bf0 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => sig00000c86,
      Q => sig00000bec
    );
  blk00000bf1 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => sig00000c85,
      Q => sig00000beb
    );
  blk00000bf2 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => sig00000c84,
      Q => sig00000bea
    );
  blk00000bf3 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => sig00000c83,
      Q => sig00000be9
    );
  blk00000bf4 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => sig00000c82,
      Q => sig00000be8
    );
  blk00000bf5 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => sig00000c81,
      Q => sig00000be7
    );
  blk00000bf6 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => sig00000c80,
      Q => sig00000be6
    );
  blk00000bf7 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => sig00000c7f,
      Q => sig00000be5
    );
  blk00000bf8 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => sig00000c7e,
      Q => sig00000c00
    );
  blk00000bf9 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => sig00000c7d,
      Q => sig00000bff
    );
  blk00000bfa : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => sig00000c7c,
      Q => sig00000bfe
    );
  blk00000bfb : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => sig00000c7b,
      Q => sig00000bfd
    );
  blk00000bfc : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => sig00000c7a,
      Q => sig00000bfc
    );
  blk00000bfd : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => sig00000c79,
      Q => sig00000bfb
    );
  blk00000bfe : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => sig00000c78,
      Q => sig00000bfa
    );
  blk00000bff : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => sig00000c77,
      Q => sig00000bf9
    );
  blk00000c00 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => sig00000c76,
      Q => sig00000bf8
    );
  blk00000c01 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => sig00000c75,
      Q => sig00000bf7
    );
  blk00000c02 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => sig00000c74,
      Q => sig00000bf6
    );
  blk00000c03 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => sig00000c73,
      Q => sig00000bf5
    );
  blk00000c04 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => sig00000c72,
      Q => sig00000bf4
    );
  blk00000c05 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => sig00000c71,
      Q => sig00000bf3
    );
  blk00000c97 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => sig00000a38,
      Q => sig00000ca0
    );
  blk00000c98 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => sig00000a37,
      Q => sig00000c9f
    );
  blk00000c99 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => sig00000a3a,
      Q => sig00000ca2
    );
  blk00000c9a : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => sig00000a39,
      Q => sig00000ca1
    );
  blk00000cab : LUT6
    generic map(
      INIT => X"FF00F0F0CCCCAAAA"
    )
    port map (
      I0 => sig000008b6,
      I1 => sig000008b6,
      I2 => sig00000ca1,
      I3 => sig00000c9b,
      I4 => sig00000c9f,
      I5 => sig00000ca0,
      O => sig00000ca3
    );
  blk00000cac : LUT6
    generic map(
      INIT => X"FF00F0F0CCCCAAAA"
    )
    port map (
      I0 => sig000008b6,
      I1 => sig00000ca1,
      I2 => sig00000ca2,
      I3 => sig00000c9c,
      I4 => sig00000c9f,
      I5 => sig00000ca0,
      O => sig00000ca4
    );
  blk00000cad : LUT6
    generic map(
      INIT => X"FF00F0F0CCCCAAAA"
    )
    port map (
      I0 => sig000008b6,
      I1 => sig00000ca2,
      I2 => sig000008b6,
      I3 => sig00000c9d,
      I4 => sig00000c9f,
      I5 => sig00000ca0,
      O => sig00000ca5
    );
  blk00000cae : LUT6
    generic map(
      INIT => X"FF00F0F0CCCCAAAA"
    )
    port map (
      I0 => sig000008b6,
      I1 => sig000008b6,
      I2 => sig000008b6,
      I3 => sig00000c9e,
      I4 => sig00000c9f,
      I5 => sig00000ca0,
      O => sig00000ca6
    );
  blk00000caf : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => sig00000ca3,
      R => sig000008b6,
      Q => sig00000c98
    );
  blk00000cb0 : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => sig00000ca4,
      R => sig000008b6,
      Q => sig00000c99
    );
  blk00000cb1 : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => sig00000ca5,
      R => sig000008b6,
      Q => sig00000c9a
    );
  blk00000cb2 : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => sig00000ca6,
      R => sig000008b6,
      Q => sig00000c97
    );
  blk00000cec : FDR
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      D => sig00000ca8,
      R => sig000008b6,
      Q => sig000000aa
    );
  blk00000ced : FD
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      D => sig00000ca9,
      Q => sig00000cc9
    );
  blk00000d5d : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => sig00000cfb,
      R => sig000008b6,
      Q => sig00000d21
    );
  blk00000d5e : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => sig00000cfa,
      R => sig000008b6,
      Q => sig00000d22
    );
  blk00000d5f : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => sig00000cf9,
      R => sig000008b6,
      Q => sig00000d23
    );
  blk00000d60 : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => sig00000cf8,
      R => sig000008b6,
      Q => sig00000d24
    );
  blk00000d61 : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => sig00000cf7,
      R => sig000008b6,
      Q => sig00000d25
    );
  blk00000d62 : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => sig00000cf6,
      R => sig000008b6,
      Q => sig00000d26
    );
  blk00000d63 : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => sig00000cf5,
      R => sig000008b6,
      Q => sig00000d27
    );
  blk00000d64 : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => sig00000cf4,
      R => sig000008b6,
      Q => sig00000d28
    );
  blk00000d65 : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => sig00000cf3,
      R => sig000008b6,
      Q => sig00000d29
    );
  blk00000d66 : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => sig00000cf2,
      R => sig000008b6,
      Q => sig00000d2a
    );
  blk00000d67 : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => sig00000cf1,
      R => sig000008b6,
      Q => sig00000d2b
    );
  blk00000d68 : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => sig00000cf0,
      R => sig000008b6,
      Q => sig00000d2c
    );
  blk00000d69 : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => sig00000cef,
      R => sig000008b6,
      Q => sig00000d2d
    );
  blk00000d6a : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => sig00000d08,
      R => sig000008b6,
      Q => sig00000cd5
    );
  blk00000d6b : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => sig00000d07,
      R => sig000008b6,
      Q => sig00000cd6
    );
  blk00000d6c : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => sig00000d06,
      R => sig000008b6,
      Q => sig00000cd7
    );
  blk00000d6d : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => sig00000d05,
      R => sig000008b6,
      Q => sig00000cd8
    );
  blk00000d6e : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => sig00000d04,
      R => sig000008b6,
      Q => sig00000cd9
    );
  blk00000d6f : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => sig00000d03,
      R => sig000008b6,
      Q => sig00000cda
    );
  blk00000d70 : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => sig00000d02,
      R => sig000008b6,
      Q => sig00000cdb
    );
  blk00000d71 : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => sig00000d01,
      R => sig000008b6,
      Q => sig00000cdc
    );
  blk00000d72 : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => sig00000d00,
      R => sig000008b6,
      Q => sig00000cdd
    );
  blk00000d73 : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => sig00000cff,
      R => sig000008b6,
      Q => sig00000cde
    );
  blk00000d74 : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => sig00000cfe,
      R => sig000008b6,
      Q => sig00000cdf
    );
  blk00000d75 : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => sig00000cfd,
      R => sig000008b6,
      Q => sig00000ce0
    );
  blk00000d76 : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => sig00000cfc,
      R => sig000008b6,
      Q => sig00000ce1
    );
  blk00000d77 : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => sig00000d14,
      R => sig000008b6,
      Q => sig00000d7c
    );
  blk00000d78 : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => sig00000d13,
      R => sig000008b6,
      Q => sig00000d7d
    );
  blk00000d79 : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => sig00000d12,
      R => sig000008b6,
      Q => sig00000d7e
    );
  blk00000d7a : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => sig00000d11,
      R => sig000008b6,
      Q => sig00000d7f
    );
  blk00000d7b : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => sig00000d10,
      R => sig000008b6,
      Q => sig00000d80
    );
  blk00000d7c : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => sig00000d0f,
      R => sig000008b6,
      Q => sig00000d81
    );
  blk00000d7d : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => sig00000d0e,
      R => sig000008b6,
      Q => sig00000d82
    );
  blk00000d7e : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => sig00000d0d,
      R => sig000008b6,
      Q => sig00000d83
    );
  blk00000d7f : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => sig00000d0c,
      R => sig000008b6,
      Q => sig00000d84
    );
  blk00000d80 : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => sig00000d0b,
      R => sig000008b6,
      Q => sig00000d85
    );
  blk00000d81 : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => sig00000d0a,
      R => sig000008b6,
      Q => sig00000d86
    );
  blk00000d82 : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => sig00000d09,
      R => sig000008b6,
      Q => sig00000d87
    );
  blk00000d83 : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => sig00000d20,
      R => sig000008b6,
      Q => sig00000d70
    );
  blk00000d84 : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => sig00000d1f,
      R => sig000008b6,
      Q => sig00000d71
    );
  blk00000d85 : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => sig00000d1e,
      R => sig000008b6,
      Q => sig00000d72
    );
  blk00000d86 : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => sig00000d1d,
      R => sig000008b6,
      Q => sig00000d73
    );
  blk00000d87 : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => sig00000d1c,
      R => sig000008b6,
      Q => sig00000d74
    );
  blk00000d88 : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => sig00000d1b,
      R => sig000008b6,
      Q => sig00000d75
    );
  blk00000d89 : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => sig00000d1a,
      R => sig000008b6,
      Q => sig00000d76
    );
  blk00000d8a : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => sig00000d19,
      R => sig000008b6,
      Q => sig00000d77
    );
  blk00000d8b : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => sig00000d18,
      R => sig000008b6,
      Q => sig00000d78
    );
  blk00000d8c : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => sig00000d17,
      R => sig000008b6,
      Q => sig00000d79
    );
  blk00000d8d : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => sig00000d16,
      R => sig000008b6,
      Q => sig00000d7a
    );
  blk00000d8e : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => sig00000d15,
      R => sig000008b6,
      Q => sig00000d7b
    );
  blk00000d8f : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => sig00000d63,
      Q => sig00000d62
    );
  blk00000d90 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => sig000000ec,
      Q => sig00000d63
    );
  blk00000eb1 : MUXCY
    port map (
      CI => sig00000de9,
      DI => sig000008b6,
      S => sig00000dc0,
      O => sig00000dce
    );
  blk00000eb2 : XORCY
    port map (
      CI => sig00000de9,
      LI => sig00000dc0,
      O => sig00000dcf
    );
  blk00000eb3 : MUXCY
    port map (
      CI => sig00000dce,
      DI => sig000008b6,
      S => sig00000dc1,
      O => sig00000dd0
    );
  blk00000eb4 : XORCY
    port map (
      CI => sig00000dce,
      LI => sig00000dc1,
      O => sig00000dd1
    );
  blk00000eb5 : MUXCY
    port map (
      CI => sig00000dd0,
      DI => sig000008b6,
      S => sig00000dc2,
      O => sig00000dd2
    );
  blk00000eb6 : XORCY
    port map (
      CI => sig00000dd0,
      LI => sig00000dc2,
      O => sig00000dd3
    );
  blk00000eb7 : MUXCY
    port map (
      CI => sig00000dd2,
      DI => sig000008b6,
      S => sig00000dc3,
      O => sig00000dd4
    );
  blk00000eb8 : XORCY
    port map (
      CI => sig00000dd2,
      LI => sig00000dc3,
      O => sig00000dd5
    );
  blk00000eb9 : MUXCY
    port map (
      CI => sig00000dd4,
      DI => sig000008b6,
      S => sig00000dc4,
      O => sig00000dd6
    );
  blk00000eba : XORCY
    port map (
      CI => sig00000dd4,
      LI => sig00000dc4,
      O => sig00000dd7
    );
  blk00000ebb : MUXCY
    port map (
      CI => sig00000dd6,
      DI => sig000008b6,
      S => sig00000dc5,
      O => sig00000dd8
    );
  blk00000ebc : XORCY
    port map (
      CI => sig00000dd6,
      LI => sig00000dc5,
      O => sig00000dd9
    );
  blk00000ebd : MUXCY
    port map (
      CI => sig00000dd8,
      DI => sig000008b6,
      S => sig00000dc6,
      O => sig00000dda
    );
  blk00000ebe : XORCY
    port map (
      CI => sig00000dd8,
      LI => sig00000dc6,
      O => sig00000ddb
    );
  blk00000ebf : MUXCY
    port map (
      CI => sig00000dda,
      DI => sig000008b6,
      S => sig00000dc7,
      O => sig00000ddc
    );
  blk00000ec0 : XORCY
    port map (
      CI => sig00000dda,
      LI => sig00000dc7,
      O => sig00000ddd
    );
  blk00000ec1 : MUXCY
    port map (
      CI => sig00000ddc,
      DI => sig000008b6,
      S => sig00000dc8,
      O => sig00000dde
    );
  blk00000ec2 : XORCY
    port map (
      CI => sig00000ddc,
      LI => sig00000dc8,
      O => sig00000ddf
    );
  blk00000ec3 : MUXCY
    port map (
      CI => sig00000dde,
      DI => sig000008b6,
      S => sig00000dc9,
      O => sig00000de0
    );
  blk00000ec4 : XORCY
    port map (
      CI => sig00000dde,
      LI => sig00000dc9,
      O => sig00000de1
    );
  blk00000ec5 : MUXCY
    port map (
      CI => sig00000de0,
      DI => sig000008b6,
      S => sig00000dca,
      O => sig00000de2
    );
  blk00000ec6 : XORCY
    port map (
      CI => sig00000de0,
      LI => sig00000dca,
      O => sig00000de3
    );
  blk00000ec7 : MUXCY
    port map (
      CI => sig00000de2,
      DI => sig000008b6,
      S => sig00000dcb,
      O => sig00000de4
    );
  blk00000ec8 : XORCY
    port map (
      CI => sig00000de2,
      LI => sig00000dcb,
      O => sig00000de5
    );
  blk00000ec9 : MUXCY
    port map (
      CI => sig00000de4,
      DI => sig000008b6,
      S => sig00000ef5,
      O => sig00000de6
    );
  blk00000eca : XORCY
    port map (
      CI => sig00000de4,
      LI => sig00000ef5,
      O => sig00000de7
    );
  blk00000ecb : MUXCY
    port map (
      CI => sig00000de6,
      DI => sig000008b6,
      S => sig00000dcc,
      O => NLW_blk00000ecb_O_UNCONNECTED
    );
  blk00000ecc : XORCY
    port map (
      CI => sig00000de6,
      LI => sig00000dcc,
      O => sig00000de8
    );
  blk00000ecd : MUXCY
    port map (
      CI => sig000006d1,
      DI => sig000008b6,
      S => sig00000dcd,
      O => sig00000de9
    );
  blk00000ece : MUXCY
    port map (
      CI => sig00000e13,
      DI => sig000008b6,
      S => sig00000dea,
      O => sig00000df8
    );
  blk00000ecf : XORCY
    port map (
      CI => sig00000e13,
      LI => sig00000dea,
      O => sig00000df9
    );
  blk00000ed0 : MUXCY
    port map (
      CI => sig00000df8,
      DI => sig000008b6,
      S => sig00000deb,
      O => sig00000dfa
    );
  blk00000ed1 : XORCY
    port map (
      CI => sig00000df8,
      LI => sig00000deb,
      O => sig00000dfb
    );
  blk00000ed2 : MUXCY
    port map (
      CI => sig00000dfa,
      DI => sig000008b6,
      S => sig00000dec,
      O => sig00000dfc
    );
  blk00000ed3 : XORCY
    port map (
      CI => sig00000dfa,
      LI => sig00000dec,
      O => sig00000dfd
    );
  blk00000ed4 : MUXCY
    port map (
      CI => sig00000dfc,
      DI => sig000008b6,
      S => sig00000ded,
      O => sig00000dfe
    );
  blk00000ed5 : XORCY
    port map (
      CI => sig00000dfc,
      LI => sig00000ded,
      O => sig00000dff
    );
  blk00000ed6 : MUXCY
    port map (
      CI => sig00000dfe,
      DI => sig000008b6,
      S => sig00000dee,
      O => sig00000e00
    );
  blk00000ed7 : XORCY
    port map (
      CI => sig00000dfe,
      LI => sig00000dee,
      O => sig00000e01
    );
  blk00000ed8 : MUXCY
    port map (
      CI => sig00000e00,
      DI => sig000008b6,
      S => sig00000def,
      O => sig00000e02
    );
  blk00000ed9 : XORCY
    port map (
      CI => sig00000e00,
      LI => sig00000def,
      O => sig00000e03
    );
  blk00000eda : MUXCY
    port map (
      CI => sig00000e02,
      DI => sig000008b6,
      S => sig00000df0,
      O => sig00000e04
    );
  blk00000edb : XORCY
    port map (
      CI => sig00000e02,
      LI => sig00000df0,
      O => sig00000e05
    );
  blk00000edc : MUXCY
    port map (
      CI => sig00000e04,
      DI => sig000008b6,
      S => sig00000df1,
      O => sig00000e06
    );
  blk00000edd : XORCY
    port map (
      CI => sig00000e04,
      LI => sig00000df1,
      O => sig00000e07
    );
  blk00000ede : MUXCY
    port map (
      CI => sig00000e06,
      DI => sig000008b6,
      S => sig00000df2,
      O => sig00000e08
    );
  blk00000edf : XORCY
    port map (
      CI => sig00000e06,
      LI => sig00000df2,
      O => sig00000e09
    );
  blk00000ee0 : MUXCY
    port map (
      CI => sig00000e08,
      DI => sig000008b6,
      S => sig00000df3,
      O => sig00000e0a
    );
  blk00000ee1 : XORCY
    port map (
      CI => sig00000e08,
      LI => sig00000df3,
      O => sig00000e0b
    );
  blk00000ee2 : MUXCY
    port map (
      CI => sig00000e0a,
      DI => sig000008b6,
      S => sig00000df4,
      O => sig00000e0c
    );
  blk00000ee3 : XORCY
    port map (
      CI => sig00000e0a,
      LI => sig00000df4,
      O => sig00000e0d
    );
  blk00000ee4 : MUXCY
    port map (
      CI => sig00000e0c,
      DI => sig000008b6,
      S => sig00000df5,
      O => sig00000e0e
    );
  blk00000ee5 : XORCY
    port map (
      CI => sig00000e0c,
      LI => sig00000df5,
      O => sig00000e0f
    );
  blk00000ee6 : MUXCY
    port map (
      CI => sig00000e0e,
      DI => sig000008b6,
      S => sig00000ef6,
      O => sig00000e10
    );
  blk00000ee7 : XORCY
    port map (
      CI => sig00000e0e,
      LI => sig00000ef6,
      O => sig00000e11
    );
  blk00000ee8 : MUXCY
    port map (
      CI => sig00000e10,
      DI => sig000008b6,
      S => sig00000df6,
      O => NLW_blk00000ee8_O_UNCONNECTED
    );
  blk00000ee9 : XORCY
    port map (
      CI => sig00000e10,
      LI => sig00000df6,
      O => sig00000e12
    );
  blk00000eea : MUXCY
    port map (
      CI => sig000006d1,
      DI => sig000008b6,
      S => sig00000df7,
      O => sig00000e13
    );
  blk00000eeb : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => sig00000d95,
      R => sig000008b6,
      Q => sig00000e69
    );
  blk00000eec : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => sig00000d94,
      R => sig000008b6,
      Q => sig00000e6a
    );
  blk00000eed : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => sig00000d93,
      R => sig000008b6,
      Q => sig00000e6b
    );
  blk00000eee : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => sig00000d92,
      R => sig000008b6,
      Q => sig00000e6c
    );
  blk00000eef : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => sig00000d91,
      R => sig000008b6,
      Q => sig00000e6d
    );
  blk00000ef0 : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => sig00000d90,
      R => sig000008b6,
      Q => sig00000e6e
    );
  blk00000ef1 : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => sig00000d8f,
      R => sig000008b6,
      Q => sig00000e6f
    );
  blk00000ef2 : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => sig00000d8e,
      R => sig000008b6,
      Q => sig00000e70
    );
  blk00000ef3 : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => sig00000d8d,
      R => sig000008b6,
      Q => sig00000e71
    );
  blk00000ef4 : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => sig00000d8c,
      R => sig000008b6,
      Q => sig00000e72
    );
  blk00000ef5 : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => sig00000d8b,
      R => sig000008b6,
      Q => sig00000e73
    );
  blk00000ef6 : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => sig00000d8a,
      R => sig000008b6,
      Q => sig00000e74
    );
  blk00000ef7 : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => sig00000d89,
      R => sig000008b6,
      Q => sig00000e75
    );
  blk00000ef8 : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => sig00000d88,
      R => sig000008b6,
      Q => sig00000e76
    );
  blk00000ef9 : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => sig00000da3,
      R => sig000008b6,
      Q => sig00000e5b
    );
  blk00000efa : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => sig00000da2,
      R => sig000008b6,
      Q => sig00000e5c
    );
  blk00000efb : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => sig00000da1,
      R => sig000008b6,
      Q => sig00000e5d
    );
  blk00000efc : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => sig00000da0,
      R => sig000008b6,
      Q => sig00000e5e
    );
  blk00000efd : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => sig00000d9f,
      R => sig000008b6,
      Q => sig00000e5f
    );
  blk00000efe : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => sig00000d9e,
      R => sig000008b6,
      Q => sig00000e60
    );
  blk00000eff : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => sig00000d9d,
      R => sig000008b6,
      Q => sig00000e61
    );
  blk00000f00 : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => sig00000d9c,
      R => sig000008b6,
      Q => sig00000e62
    );
  blk00000f01 : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => sig00000d9b,
      R => sig000008b6,
      Q => sig00000e63
    );
  blk00000f02 : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => sig00000d9a,
      R => sig000008b6,
      Q => sig00000e64
    );
  blk00000f03 : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => sig00000d99,
      R => sig000008b6,
      Q => sig00000e65
    );
  blk00000f04 : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => sig00000d98,
      R => sig000008b6,
      Q => sig00000e66
    );
  blk00000f05 : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => sig00000d97,
      R => sig000008b6,
      Q => sig00000e67
    );
  blk00000f06 : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => sig00000d96,
      R => sig000008b6,
      Q => sig00000e68
    );
  blk00000f07 : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => sig00000db1,
      R => sig000008b6,
      Q => sig00000e23
    );
  blk00000f08 : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => sig00000db0,
      R => sig000008b6,
      Q => sig00000e24
    );
  blk00000f09 : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => sig00000daf,
      R => sig000008b6,
      Q => sig00000e25
    );
  blk00000f0a : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => sig00000dae,
      R => sig000008b6,
      Q => sig00000e26
    );
  blk00000f0b : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => sig00000dad,
      R => sig000008b6,
      Q => sig00000e27
    );
  blk00000f0c : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => sig00000dac,
      R => sig000008b6,
      Q => sig00000e28
    );
  blk00000f0d : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => sig00000dab,
      R => sig000008b6,
      Q => sig00000e29
    );
  blk00000f0e : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => sig00000daa,
      R => sig000008b6,
      Q => sig00000e2a
    );
  blk00000f0f : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => sig00000da9,
      R => sig000008b6,
      Q => sig00000e2b
    );
  blk00000f10 : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => sig00000da8,
      R => sig000008b6,
      Q => sig00000e2c
    );
  blk00000f11 : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => sig00000da7,
      R => sig000008b6,
      Q => sig00000e2d
    );
  blk00000f12 : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => sig00000da6,
      R => sig000008b6,
      Q => sig00000e2e
    );
  blk00000f13 : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => sig00000da5,
      R => sig000008b6,
      Q => sig00000e2f
    );
  blk00000f14 : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => sig00000da4,
      R => sig000008b6,
      Q => sig00000e30
    );
  blk00000f15 : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => sig00000dbf,
      R => sig000008b6,
      Q => sig00000caa
    );
  blk00000f16 : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => sig00000dbe,
      R => sig000008b6,
      Q => sig00000cab
    );
  blk00000f17 : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => sig00000dbd,
      R => sig000008b6,
      Q => sig00000cac
    );
  blk00000f18 : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => sig00000dbc,
      R => sig000008b6,
      Q => sig00000cad
    );
  blk00000f19 : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => sig00000dbb,
      R => sig000008b6,
      Q => sig00000cae
    );
  blk00000f1a : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => sig00000dba,
      R => sig000008b6,
      Q => sig00000caf
    );
  blk00000f1b : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => sig00000db9,
      R => sig000008b6,
      Q => sig00000cb0
    );
  blk00000f1c : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => sig00000db8,
      R => sig000008b6,
      Q => sig00000cb1
    );
  blk00000f1d : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => sig00000db7,
      R => sig000008b6,
      Q => sig00000cb2
    );
  blk00000f1e : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => sig00000db6,
      R => sig000008b6,
      Q => sig00000cb3
    );
  blk00000f1f : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => sig00000db5,
      R => sig000008b6,
      Q => sig00000cb4
    );
  blk00000f20 : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => sig00000db4,
      R => sig000008b6,
      Q => sig00000cb5
    );
  blk00000f21 : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => sig00000db3,
      R => sig000008b6,
      Q => sig00000cb6
    );
  blk00000f22 : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => sig00000db2,
      R => sig000008b6,
      Q => sig00000cb7
    );
  blk00000f23 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => sig00000dcf,
      Q => sig00000e93
    );
  blk00000f24 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => sig00000dd1,
      Q => sig00000e94
    );
  blk00000f25 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => sig00000dd3,
      Q => sig00000e95
    );
  blk00000f26 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => sig00000dd5,
      Q => sig00000e96
    );
  blk00000f27 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => sig00000dd7,
      Q => sig00000e97
    );
  blk00000f28 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => sig00000dd9,
      Q => sig00000e98
    );
  blk00000f29 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => sig00000ddb,
      Q => sig00000e99
    );
  blk00000f2a : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => sig00000ddd,
      Q => sig00000e9a
    );
  blk00000f2b : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => sig00000ddf,
      Q => sig00000e9b
    );
  blk00000f2c : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => sig00000de1,
      Q => sig00000e9c
    );
  blk00000f2d : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => sig00000de3,
      Q => sig00000e9d
    );
  blk00000f2e : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => sig00000de5,
      Q => sig00000e9e
    );
  blk00000f2f : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => sig00000de7,
      Q => sig00000e9f
    );
  blk00000f30 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => sig00000de8,
      Q => sig00000ea0
    );
  blk00000f31 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => sig00000df9,
      Q => sig00000ea1
    );
  blk00000f32 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => sig00000dfb,
      Q => sig00000ea2
    );
  blk00000f33 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => sig00000dfd,
      Q => sig00000ea3
    );
  blk00000f34 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => sig00000dff,
      Q => sig00000ea4
    );
  blk00000f35 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => sig00000e01,
      Q => sig00000ea5
    );
  blk00000f36 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => sig00000e03,
      Q => sig00000ea6
    );
  blk00000f37 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => sig00000e05,
      Q => sig00000ea7
    );
  blk00000f38 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => sig00000e07,
      Q => sig00000ea8
    );
  blk00000f39 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => sig00000e09,
      Q => sig00000ea9
    );
  blk00000f3a : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => sig00000e0b,
      Q => sig00000eaa
    );
  blk00000f3b : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => sig00000e0d,
      Q => sig00000eab
    );
  blk00000f3c : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => sig00000e0f,
      Q => sig00000eac
    );
  blk00000f3d : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => sig00000e11,
      Q => sig00000ead
    );
  blk00000f3e : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => sig00000e12,
      Q => sig00000eae
    );
  blk00000f3f : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => sig00000cc8,
      Q => sig00000eb4
    );
  blk00000f40 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => sig00000eb1,
      Q => sig00000eb0
    );
  blk00000f41 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => sig00000e14,
      Q => sig00000eaf
    );
  blk00000f42 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => sig00000cd3,
      Q => sig00000eb3
    );
  blk00000f43 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => sig00000eae,
      Q => sig00000e22
    );
  blk00000f44 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => sig00000ead,
      Q => sig00000e21
    );
  blk00000f45 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => sig00000eac,
      Q => sig00000e20
    );
  blk00000f46 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => sig00000eab,
      Q => sig00000e1f
    );
  blk00000f47 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => sig00000eaa,
      Q => sig00000e1e
    );
  blk00000f48 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => sig00000ea9,
      Q => sig00000e1d
    );
  blk00000f49 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => sig00000ea8,
      Q => sig00000e1c
    );
  blk00000f4a : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => sig00000ea7,
      Q => sig00000e1b
    );
  blk00000f4b : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => sig00000ea6,
      Q => sig00000e1a
    );
  blk00000f4c : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => sig00000ea5,
      Q => sig00000e19
    );
  blk00000f4d : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => sig00000ea4,
      Q => sig00000e18
    );
  blk00000f4e : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => sig00000ea3,
      Q => sig00000e17
    );
  blk00000f4f : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => sig00000ea2,
      Q => sig00000e16
    );
  blk00000f50 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => sig00000ea1,
      Q => sig00000e15
    );
  blk00000f51 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => sig00000e30,
      Q => sig00000cc5
    );
  blk00000f52 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => sig00000e2f,
      Q => sig00000cc4
    );
  blk00000f53 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => sig00000e2e,
      Q => sig00000cc3
    );
  blk00000f54 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => sig00000e2d,
      Q => sig00000cc2
    );
  blk00000f55 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => sig00000e2c,
      Q => sig00000cc1
    );
  blk00000f56 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => sig00000e2b,
      Q => sig00000cc0
    );
  blk00000f57 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => sig00000e2a,
      Q => sig00000cbf
    );
  blk00000f58 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => sig00000e29,
      Q => sig00000cbe
    );
  blk00000f59 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => sig00000e28,
      Q => sig00000cbd
    );
  blk00000f5a : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => sig00000e27,
      Q => sig00000cbc
    );
  blk00000f5b : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => sig00000e26,
      Q => sig00000cbb
    );
  blk00000f5c : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => sig00000e25,
      Q => sig00000cba
    );
  blk00000f5d : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => sig00000e24,
      Q => sig00000cb9
    );
  blk00000f5e : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => sig00000e23,
      Q => sig00000cb8
    );
  blk00000f5f : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => sig00000e4c,
      Q => sig00000e3e
    );
  blk00000f60 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => sig00000e4b,
      Q => sig00000e3d
    );
  blk00000f61 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => sig00000e4a,
      Q => sig00000e3c
    );
  blk00000f62 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => sig00000e49,
      Q => sig00000e3b
    );
  blk00000f63 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => sig00000e48,
      Q => sig00000e3a
    );
  blk00000f64 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => sig00000e47,
      Q => sig00000e39
    );
  blk00000f65 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => sig00000e46,
      Q => sig00000e38
    );
  blk00000f66 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => sig00000e45,
      Q => sig00000e37
    );
  blk00000f67 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => sig00000e44,
      Q => sig00000e36
    );
  blk00000f68 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => sig00000e43,
      Q => sig00000e35
    );
  blk00000f69 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => sig00000e42,
      Q => sig00000e34
    );
  blk00000f6a : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => sig00000e41,
      Q => sig00000e33
    );
  blk00000f6b : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => sig00000e40,
      Q => sig00000e32
    );
  blk00000f6c : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => sig00000e3f,
      Q => sig00000e31
    );
  blk00000f6d : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => sig00000e76,
      Q => sig00000e92
    );
  blk00000f6e : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => sig00000e75,
      Q => sig00000e91
    );
  blk00000f6f : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => sig00000e74,
      Q => sig00000e90
    );
  blk00000f70 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => sig00000e73,
      Q => sig00000e8f
    );
  blk00000f71 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => sig00000e72,
      Q => sig00000e8e
    );
  blk00000f72 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => sig00000e71,
      Q => sig00000e8d
    );
  blk00000f73 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => sig00000e70,
      Q => sig00000e8c
    );
  blk00000f74 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => sig00000e6f,
      Q => sig00000e8b
    );
  blk00000f75 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => sig00000e6e,
      Q => sig00000e8a
    );
  blk00000f76 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => sig00000e6d,
      Q => sig00000e89
    );
  blk00000f77 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => sig00000e6c,
      Q => sig00000e88
    );
  blk00000f78 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => sig00000e6b,
      Q => sig00000e87
    );
  blk00000f79 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => sig00000e6a,
      Q => sig00000e86
    );
  blk00000f7a : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => sig00000e69,
      Q => sig00000e85
    );
  blk00000f7b : LUT6
    generic map(
      INIT => X"FF00F0F0CCCCAAAA"
    )
    port map (
      I0 => sig000008b6,
      I1 => sig000008b6,
      I2 => sig000008b6,
      I3 => sig00000cb8,
      I4 => sig00000cc6,
      I5 => sig00000cc7,
      O => sig00000eb5
    );
  blk00000f7c : LUT6
    generic map(
      INIT => X"FF00F0F0CCCCAAAA"
    )
    port map (
      I0 => sig000008b6,
      I1 => sig000008b6,
      I2 => sig00000cb8,
      I3 => sig00000cb9,
      I4 => sig00000cc6,
      I5 => sig00000cc7,
      O => sig00000eb6
    );
  blk00000f7d : LUT6
    generic map(
      INIT => X"FF00F0F0CCCCAAAA"
    )
    port map (
      I0 => sig000008b6,
      I1 => sig00000cb8,
      I2 => sig00000cb9,
      I3 => sig00000cba,
      I4 => sig00000cc6,
      I5 => sig00000cc7,
      O => sig00000eb7
    );
  blk00000f7e : LUT6
    generic map(
      INIT => X"FF00F0F0CCCCAAAA"
    )
    port map (
      I0 => sig00000cb8,
      I1 => sig00000cb9,
      I2 => sig00000cba,
      I3 => sig00000cbb,
      I4 => sig00000cc6,
      I5 => sig00000cc7,
      O => sig00000eb8
    );
  blk00000f7f : LUT6
    generic map(
      INIT => X"FF00F0F0CCCCAAAA"
    )
    port map (
      I0 => sig00000cb9,
      I1 => sig00000cba,
      I2 => sig00000cbb,
      I3 => sig00000cbc,
      I4 => sig00000cc6,
      I5 => sig00000cc7,
      O => sig00000eb9
    );
  blk00000f80 : LUT6
    generic map(
      INIT => X"FF00F0F0CCCCAAAA"
    )
    port map (
      I0 => sig00000cba,
      I1 => sig00000cbb,
      I2 => sig00000cbc,
      I3 => sig00000cbd,
      I4 => sig00000cc6,
      I5 => sig00000cc7,
      O => sig00000eba
    );
  blk00000f81 : LUT6
    generic map(
      INIT => X"FF00F0F0CCCCAAAA"
    )
    port map (
      I0 => sig00000cbb,
      I1 => sig00000cbc,
      I2 => sig00000cbd,
      I3 => sig00000cbe,
      I4 => sig00000cc6,
      I5 => sig00000cc7,
      O => sig00000ebb
    );
  blk00000f82 : LUT6
    generic map(
      INIT => X"FF00F0F0CCCCAAAA"
    )
    port map (
      I0 => sig00000cbc,
      I1 => sig00000cbd,
      I2 => sig00000cbe,
      I3 => sig00000cbf,
      I4 => sig00000cc6,
      I5 => sig00000cc7,
      O => sig00000ebc
    );
  blk00000f83 : LUT6
    generic map(
      INIT => X"FF00F0F0CCCCAAAA"
    )
    port map (
      I0 => sig00000cbd,
      I1 => sig00000cbe,
      I2 => sig00000cbf,
      I3 => sig00000cc0,
      I4 => sig00000cc6,
      I5 => sig00000cc7,
      O => sig00000ebd
    );
  blk00000f84 : LUT6
    generic map(
      INIT => X"FF00F0F0CCCCAAAA"
    )
    port map (
      I0 => sig00000cbe,
      I1 => sig00000cbf,
      I2 => sig00000cc0,
      I3 => sig00000cc1,
      I4 => sig00000cc6,
      I5 => sig00000cc7,
      O => sig00000ebe
    );
  blk00000f85 : LUT6
    generic map(
      INIT => X"FF00F0F0CCCCAAAA"
    )
    port map (
      I0 => sig00000cbf,
      I1 => sig00000cc0,
      I2 => sig00000cc1,
      I3 => sig00000cc2,
      I4 => sig00000cc6,
      I5 => sig00000cc7,
      O => sig00000ebf
    );
  blk00000f86 : LUT6
    generic map(
      INIT => X"FF00F0F0CCCCAAAA"
    )
    port map (
      I0 => sig00000cc0,
      I1 => sig00000cc1,
      I2 => sig00000cc2,
      I3 => sig00000cc3,
      I4 => sig00000cc6,
      I5 => sig00000cc7,
      O => sig00000ec0
    );
  blk00000f87 : LUT6
    generic map(
      INIT => X"FF00F0F0CCCCAAAA"
    )
    port map (
      I0 => sig00000cc1,
      I1 => sig00000cc2,
      I2 => sig00000cc3,
      I3 => sig00000cc4,
      I4 => sig00000cc6,
      I5 => sig00000cc7,
      O => sig00000ec1
    );
  blk00000f88 : LUT6
    generic map(
      INIT => X"FF00F0F0CCCCAAAA"
    )
    port map (
      I0 => sig00000cc2,
      I1 => sig00000cc3,
      I2 => sig00000cc4,
      I3 => sig00000cc5,
      I4 => sig00000cc6,
      I5 => sig00000cc7,
      O => sig00000ec2
    );
  blk00000f89 : LUT6
    generic map(
      INIT => X"FF00F0F0CCCCAAAA"
    )
    port map (
      I0 => sig00000cc3,
      I1 => sig00000cc4,
      I2 => sig00000cc5,
      I3 => sig00000cc5,
      I4 => sig00000cc6,
      I5 => sig00000cc7,
      O => sig00000ec3
    );
  blk00000f8a : LUT6
    generic map(
      INIT => X"FF00F0F0CCCCAAAA"
    )
    port map (
      I0 => sig00000cc4,
      I1 => sig00000cc5,
      I2 => sig00000cc5,
      I3 => sig00000cc5,
      I4 => sig00000cc6,
      I5 => sig00000cc7,
      O => sig00000ec4
    );
  blk00000f8b : LUT6
    generic map(
      INIT => X"FF00F0F0CCCCAAAA"
    )
    port map (
      I0 => sig00000cc5,
      I1 => sig00000cc5,
      I2 => sig00000cc5,
      I3 => sig00000cc5,
      I4 => sig00000cc6,
      I5 => sig00000cc7,
      O => sig00000ec5
    );
  blk00000f8c : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => sig00000eb5,
      R => sig000008b6,
      Q => NLW_blk00000f8c_Q_UNCONNECTED
    );
  blk00000f8d : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => sig00000eb6,
      R => sig000008b6,
      Q => NLW_blk00000f8d_Q_UNCONNECTED
    );
  blk00000f8e : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => sig00000eb7,
      R => sig000008b6,
      Q => NLW_blk00000f8e_Q_UNCONNECTED
    );
  blk00000f8f : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => sig00000eb8,
      R => sig000008b6,
      Q => sig000000b7
    );
  blk00000f90 : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => sig00000eb9,
      R => sig000008b6,
      Q => sig000000b8
    );
  blk00000f91 : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => sig00000eba,
      R => sig000008b6,
      Q => sig000000b9
    );
  blk00000f92 : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => sig00000ebb,
      R => sig000008b6,
      Q => sig000000ba
    );
  blk00000f93 : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => sig00000ebc,
      R => sig000008b6,
      Q => sig000000bb
    );
  blk00000f94 : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => sig00000ebd,
      R => sig000008b6,
      Q => sig000000bc
    );
  blk00000f95 : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => sig00000ebe,
      R => sig000008b6,
      Q => sig000000bd
    );
  blk00000f96 : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => sig00000ebf,
      R => sig000008b6,
      Q => sig000000be
    );
  blk00000f97 : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => sig00000ec0,
      R => sig000008b6,
      Q => sig000000bf
    );
  blk00000f98 : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => sig00000ec1,
      R => sig000008b6,
      Q => sig000000c0
    );
  blk00000f99 : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => sig00000ec2,
      R => sig000008b6,
      Q => sig000000c1
    );
  blk00000f9a : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => sig00000ec3,
      R => sig000008b6,
      Q => sig000000c2
    );
  blk00000f9b : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => sig00000ec4,
      R => sig000008b6,
      Q => NLW_blk00000f9b_Q_UNCONNECTED
    );
  blk00000f9c : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => sig00000ec5,
      R => sig000008b6,
      Q => NLW_blk00000f9c_Q_UNCONNECTED
    );
  blk00000f9d : LUT6
    generic map(
      INIT => X"FF00F0F0CCCCAAAA"
    )
    port map (
      I0 => sig000008b6,
      I1 => sig000008b6,
      I2 => sig000008b6,
      I3 => sig00000caa,
      I4 => sig00000cc6,
      I5 => sig00000cc7,
      O => sig00000ec6
    );
  blk00000f9e : LUT6
    generic map(
      INIT => X"FF00F0F0CCCCAAAA"
    )
    port map (
      I0 => sig000008b6,
      I1 => sig000008b6,
      I2 => sig00000caa,
      I3 => sig00000cab,
      I4 => sig00000cc6,
      I5 => sig00000cc7,
      O => sig00000ec7
    );
  blk00000f9f : LUT6
    generic map(
      INIT => X"FF00F0F0CCCCAAAA"
    )
    port map (
      I0 => sig000008b6,
      I1 => sig00000caa,
      I2 => sig00000cab,
      I3 => sig00000cac,
      I4 => sig00000cc6,
      I5 => sig00000cc7,
      O => sig00000ec8
    );
  blk00000fa0 : LUT6
    generic map(
      INIT => X"FF00F0F0CCCCAAAA"
    )
    port map (
      I0 => sig00000caa,
      I1 => sig00000cab,
      I2 => sig00000cac,
      I3 => sig00000cad,
      I4 => sig00000cc6,
      I5 => sig00000cc7,
      O => sig00000ec9
    );
  blk00000fa1 : LUT6
    generic map(
      INIT => X"FF00F0F0CCCCAAAA"
    )
    port map (
      I0 => sig00000cab,
      I1 => sig00000cac,
      I2 => sig00000cad,
      I3 => sig00000cae,
      I4 => sig00000cc6,
      I5 => sig00000cc7,
      O => sig00000eca
    );
  blk00000fa2 : LUT6
    generic map(
      INIT => X"FF00F0F0CCCCAAAA"
    )
    port map (
      I0 => sig00000cac,
      I1 => sig00000cad,
      I2 => sig00000cae,
      I3 => sig00000caf,
      I4 => sig00000cc6,
      I5 => sig00000cc7,
      O => sig00000ecb
    );
  blk00000fa3 : LUT6
    generic map(
      INIT => X"FF00F0F0CCCCAAAA"
    )
    port map (
      I0 => sig00000cad,
      I1 => sig00000cae,
      I2 => sig00000caf,
      I3 => sig00000cb0,
      I4 => sig00000cc6,
      I5 => sig00000cc7,
      O => sig00000ecc
    );
  blk00000fa4 : LUT6
    generic map(
      INIT => X"FF00F0F0CCCCAAAA"
    )
    port map (
      I0 => sig00000cae,
      I1 => sig00000caf,
      I2 => sig00000cb0,
      I3 => sig00000cb1,
      I4 => sig00000cc6,
      I5 => sig00000cc7,
      O => sig00000ecd
    );
  blk00000fa5 : LUT6
    generic map(
      INIT => X"FF00F0F0CCCCAAAA"
    )
    port map (
      I0 => sig00000caf,
      I1 => sig00000cb0,
      I2 => sig00000cb1,
      I3 => sig00000cb2,
      I4 => sig00000cc6,
      I5 => sig00000cc7,
      O => sig00000ece
    );
  blk00000fa6 : LUT6
    generic map(
      INIT => X"FF00F0F0CCCCAAAA"
    )
    port map (
      I0 => sig00000cb0,
      I1 => sig00000cb1,
      I2 => sig00000cb2,
      I3 => sig00000cb3,
      I4 => sig00000cc6,
      I5 => sig00000cc7,
      O => sig00000ecf
    );
  blk00000fa7 : LUT6
    generic map(
      INIT => X"FF00F0F0CCCCAAAA"
    )
    port map (
      I0 => sig00000cb1,
      I1 => sig00000cb2,
      I2 => sig00000cb3,
      I3 => sig00000cb4,
      I4 => sig00000cc6,
      I5 => sig00000cc7,
      O => sig00000ed0
    );
  blk00000fa8 : LUT6
    generic map(
      INIT => X"FF00F0F0CCCCAAAA"
    )
    port map (
      I0 => sig00000cb2,
      I1 => sig00000cb3,
      I2 => sig00000cb4,
      I3 => sig00000cb5,
      I4 => sig00000cc6,
      I5 => sig00000cc7,
      O => sig00000ed1
    );
  blk00000fa9 : LUT6
    generic map(
      INIT => X"FF00F0F0CCCCAAAA"
    )
    port map (
      I0 => sig00000cb3,
      I1 => sig00000cb4,
      I2 => sig00000cb5,
      I3 => sig00000cb6,
      I4 => sig00000cc6,
      I5 => sig00000cc7,
      O => sig00000ed2
    );
  blk00000faa : LUT6
    generic map(
      INIT => X"FF00F0F0CCCCAAAA"
    )
    port map (
      I0 => sig00000cb4,
      I1 => sig00000cb5,
      I2 => sig00000cb6,
      I3 => sig00000cb7,
      I4 => sig00000cc6,
      I5 => sig00000cc7,
      O => sig00000ed3
    );
  blk00000fab : LUT6
    generic map(
      INIT => X"FF00F0F0CCCCAAAA"
    )
    port map (
      I0 => sig00000cb5,
      I1 => sig00000cb6,
      I2 => sig00000cb7,
      I3 => sig00000cb7,
      I4 => sig00000cc6,
      I5 => sig00000cc7,
      O => sig00000ed4
    );
  blk00000fac : LUT6
    generic map(
      INIT => X"FF00F0F0CCCCAAAA"
    )
    port map (
      I0 => sig00000cb6,
      I1 => sig00000cb7,
      I2 => sig00000cb7,
      I3 => sig00000cb7,
      I4 => sig00000cc6,
      I5 => sig00000cc7,
      O => sig00000ed5
    );
  blk00000fad : LUT6
    generic map(
      INIT => X"FF00F0F0CCCCAAAA"
    )
    port map (
      I0 => sig00000cb7,
      I1 => sig00000cb7,
      I2 => sig00000cb7,
      I3 => sig00000cb7,
      I4 => sig00000cc6,
      I5 => sig00000cc7,
      O => sig00000ed6
    );
  blk00000fae : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => sig00000ec6,
      R => sig000008b6,
      Q => NLW_blk00000fae_Q_UNCONNECTED
    );
  blk00000faf : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => sig00000ec7,
      R => sig000008b6,
      Q => NLW_blk00000faf_Q_UNCONNECTED
    );
  blk00000fb0 : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => sig00000ec8,
      R => sig000008b6,
      Q => NLW_blk00000fb0_Q_UNCONNECTED
    );
  blk00000fb1 : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => sig00000ec9,
      R => sig000008b6,
      Q => sig000000ab
    );
  blk00000fb2 : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => sig00000eca,
      R => sig000008b6,
      Q => sig000000ac
    );
  blk00000fb3 : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => sig00000ecb,
      R => sig000008b6,
      Q => sig000000ad
    );
  blk00000fb4 : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => sig00000ecc,
      R => sig000008b6,
      Q => sig000000ae
    );
  blk00000fb5 : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => sig00000ecd,
      R => sig000008b6,
      Q => sig000000af
    );
  blk00000fb6 : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => sig00000ece,
      R => sig000008b6,
      Q => sig000000b0
    );
  blk00000fb7 : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => sig00000ecf,
      R => sig000008b6,
      Q => sig000000b1
    );
  blk00000fb8 : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => sig00000ed0,
      R => sig000008b6,
      Q => sig000000b2
    );
  blk00000fb9 : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => sig00000ed1,
      R => sig000008b6,
      Q => sig000000b3
    );
  blk00000fba : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => sig00000ed2,
      R => sig000008b6,
      Q => sig000000b4
    );
  blk00000fbb : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => sig00000ed3,
      R => sig000008b6,
      Q => sig000000b5
    );
  blk00000fbc : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => sig00000ed4,
      R => sig000008b6,
      Q => sig000000b6
    );
  blk00000fbd : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => sig00000ed5,
      R => sig000008b6,
      Q => NLW_blk00000fbd_Q_UNCONNECTED
    );
  blk00000fbe : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => sig00000ed6,
      R => sig000008b6,
      Q => NLW_blk00000fbe_Q_UNCONNECTED
    );
  blk00000fd2 : FDR
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      D => sig00000ed7,
      R => sig000008b6,
      Q => NlwRenamedSig_OI_xk_index(0)
    );
  blk00000fd3 : FDR
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      D => sig00000ed8,
      R => sig000008b6,
      Q => NlwRenamedSig_OI_xk_index(1)
    );
  blk00000fd4 : FDR
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      D => sig00000ed9,
      R => sig000008b6,
      Q => NlwRenamedSig_OI_xk_index(2)
    );
  blk00000fd5 : FDR
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      D => sig00000eda,
      R => sig000008b6,
      Q => NlwRenamedSig_OI_xk_index(3)
    );
  blk00000fd6 : FDR
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      D => sig00000edb,
      R => sig000008b6,
      Q => NlwRenamedSig_OI_xk_index(4)
    );
  blk00000fd7 : FDR
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      D => sig00000edc,
      R => sig000008b6,
      Q => NlwRenamedSig_OI_xk_index(5)
    );
  blk00000fdd : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => sig00000ee9,
      D => sig00000ee3,
      R => sig000008b6,
      Q => sig00000eec
    );
  blk00000fde : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => sig00000ee9,
      D => sig00000ee4,
      R => sig000008b6,
      Q => sig00000eeb
    );
  blk00000fdf : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => sig00000ee9,
      D => sig00000ee5,
      R => sig000008b6,
      Q => sig00000eea
    );
  blk00000fe0 : FDR
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      D => sig00000ee7,
      R => sig000008b6,
      Q => sig00000eed
    );
  blk00000fe1 : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => sig00000ee9,
      D => sig00000ee8,
      R => sig000008b6,
      Q => U0_i_synth_non_floating_point_arch_d_xfft_inst_has_bit_reverse_busy_gen_busy_i
    );
  blk00000fe2 : LUT4
    generic map(
      INIT => X"AA20"
    )
    port map (
      I0 => ce,
      I1 => sig0000005e,
      I2 => sig00000114,
      I3 => sig000000a3,
      O => sig00000013
    );
  blk00000fe3 : LUT3
    generic map(
      INIT => X"D8"
    )
    port map (
      I0 => ce,
      I1 => sig000000a4,
      I2 => sig0000009b,
      O => sig0000000c
    );
  blk00000fe4 : LUT3
    generic map(
      INIT => X"D8"
    )
    port map (
      I0 => ce,
      I1 => sig000000a5,
      I2 => sig0000009c,
      O => sig0000000b
    );
  blk00000fe5 : LUT3
    generic map(
      INIT => X"D8"
    )
    port map (
      I0 => ce,
      I1 => sig000000a6,
      I2 => sig0000009d,
      O => sig0000000a
    );
  blk00000fe6 : LUT3
    generic map(
      INIT => X"D8"
    )
    port map (
      I0 => ce,
      I1 => sig000000a7,
      I2 => sig0000009e,
      O => sig00000009
    );
  blk00000fe7 : LUT3
    generic map(
      INIT => X"D8"
    )
    port map (
      I0 => ce,
      I1 => sig000000a8,
      I2 => sig0000009f,
      O => sig00000008
    );
  blk00000fe8 : LUT3
    generic map(
      INIT => X"D8"
    )
    port map (
      I0 => ce,
      I1 => sig000000a9,
      I2 => sig000000a0,
      O => sig00000007
    );
  blk00000fe9 : LUT3
    generic map(
      INIT => X"D8"
    )
    port map (
      I0 => ce,
      I1 => sig000000a4,
      I2 => sig00000098,
      O => sig00000012
    );
  blk00000fea : LUT3
    generic map(
      INIT => X"D8"
    )
    port map (
      I0 => ce,
      I1 => sig000000a5,
      I2 => sig00000097,
      O => sig00000011
    );
  blk00000feb : LUT3
    generic map(
      INIT => X"D8"
    )
    port map (
      I0 => ce,
      I1 => sig000000a6,
      I2 => sig00000096,
      O => sig00000010
    );
  blk00000fec : LUT3
    generic map(
      INIT => X"D8"
    )
    port map (
      I0 => ce,
      I1 => sig000000a7,
      I2 => sig00000095,
      O => sig0000000f
    );
  blk00000fed : LUT3
    generic map(
      INIT => X"D8"
    )
    port map (
      I0 => ce,
      I1 => sig000000a8,
      I2 => sig00000094,
      O => sig0000000e
    );
  blk00000fee : LUT3
    generic map(
      INIT => X"D8"
    )
    port map (
      I0 => ce,
      I1 => sig000000a9,
      I2 => sig00000093,
      O => sig0000000d
    );
  blk00000fef : LUT3
    generic map(
      INIT => X"D8"
    )
    port map (
      I0 => ce,
      I1 => sig00000001,
      I2 => sig00000061,
      O => sig00000002
    );
  blk00000ff0 : LUT3
    generic map(
      INIT => X"D8"
    )
    port map (
      I0 => ce,
      I1 => sig00000003,
      I2 => sig00000062,
      O => sig00000004
    );
  blk00000ff1 : LUT3
    generic map(
      INIT => X"D8"
    )
    port map (
      I0 => ce,
      I1 => sig00000005,
      I2 => NlwRenamedSig_OI_cpv,
      O => sig00000006
    );
  blk00000ff2 : LUT3
    generic map(
      INIT => X"D8"
    )
    port map (
      I0 => ce,
      I1 => sig00000015,
      I2 => sig00000112,
      O => sig00000016
    );
  blk00000ff3 : LUT2
    generic map(
      INIT => X"2"
    )
    port map (
      I0 => sig0000011b,
      I1 => sig00000114,
      O => sig0000001b
    );
  blk00000ff4 : LUT2
    generic map(
      INIT => X"2"
    )
    port map (
      I0 => sig0000011a,
      I1 => sig00000114,
      O => sig0000001c
    );
  blk00000ff5 : LUT2
    generic map(
      INIT => X"2"
    )
    port map (
      I0 => sig00000119,
      I1 => sig00000114,
      O => sig0000001d
    );
  blk00000ff6 : LUT2
    generic map(
      INIT => X"2"
    )
    port map (
      I0 => sig00000118,
      I1 => sig00000114,
      O => sig0000001e
    );
  blk00000ff7 : LUT2
    generic map(
      INIT => X"2"
    )
    port map (
      I0 => sig00000117,
      I1 => sig00000114,
      O => sig0000001f
    );
  blk00000ff8 : LUT2
    generic map(
      INIT => X"4"
    )
    port map (
      I0 => sig00000114,
      I1 => sig00000116,
      O => sig00000020
    );
  blk00000ff9 : LUT3
    generic map(
      INIT => X"D8"
    )
    port map (
      I0 => sig0000009a,
      I1 => sig0000004c,
      I2 => sig00000051,
      O => sig00000033
    );
  blk00000ffa : LUT3
    generic map(
      INIT => X"D8"
    )
    port map (
      I0 => sig0000009a,
      I1 => sig0000004d,
      I2 => sig00000050,
      O => sig00000034
    );
  blk00000ffb : LUT3
    generic map(
      INIT => X"D8"
    )
    port map (
      I0 => sig0000009a,
      I1 => sig0000004e,
      I2 => sig0000004f,
      O => sig00000035
    );
  blk00000ffc : LUT3
    generic map(
      INIT => X"D8"
    )
    port map (
      I0 => sig0000009a,
      I1 => sig0000004f,
      I2 => sig0000004e,
      O => sig00000036
    );
  blk00000ffd : LUT3
    generic map(
      INIT => X"D8"
    )
    port map (
      I0 => sig0000009a,
      I1 => sig00000050,
      I2 => sig0000004d,
      O => sig00000037
    );
  blk00000ffe : LUT3
    generic map(
      INIT => X"D8"
    )
    port map (
      I0 => sig0000009a,
      I1 => sig00000051,
      I2 => sig0000004c,
      O => sig00000038
    );
  blk00000fff : LUT3
    generic map(
      INIT => X"D8"
    )
    port map (
      I0 => sig00000099,
      I1 => sig0000009b,
      I2 => sig00000093,
      O => sig00000039
    );
  blk00001000 : LUT3
    generic map(
      INIT => X"D8"
    )
    port map (
      I0 => sig00000099,
      I1 => sig0000009c,
      I2 => sig00000094,
      O => sig0000003a
    );
  blk00001001 : LUT3
    generic map(
      INIT => X"D8"
    )
    port map (
      I0 => sig00000099,
      I1 => sig0000009d,
      I2 => sig00000095,
      O => sig0000003b
    );
  blk00001002 : LUT3
    generic map(
      INIT => X"D8"
    )
    port map (
      I0 => sig00000099,
      I1 => sig0000009e,
      I2 => sig00000096,
      O => sig0000003c
    );
  blk00001003 : LUT3
    generic map(
      INIT => X"D8"
    )
    port map (
      I0 => sig00000099,
      I1 => sig0000009f,
      I2 => sig00000097,
      O => sig0000003d
    );
  blk00001004 : LUT3
    generic map(
      INIT => X"D8"
    )
    port map (
      I0 => sig00000099,
      I1 => sig000000a0,
      I2 => sig00000098,
      O => sig0000003e
    );
  blk00001005 : LUT2
    generic map(
      INIT => X"8"
    )
    port map (
      I0 => sig00000115,
      I1 => ce,
      O => sig00000017
    );
  blk00001006 : LUT2
    generic map(
      INIT => X"E"
    )
    port map (
      I0 => sig00000047,
      I1 => sig00000114,
      O => sig00000042
    );
  blk00001007 : LUT2
    generic map(
      INIT => X"2"
    )
    port map (
      I0 => sig00000f16,
      I1 => sig0000005e,
      O => sig00000043
    );
  blk00001008 : LUT2
    generic map(
      INIT => X"4"
    )
    port map (
      I0 => sig00000049,
      I1 => ce,
      O => sig00000044
    );
  blk00001009 : LUT5
    generic map(
      INIT => X"B000B0B0"
    )
    port map (
      I0 => sig00000191,
      I1 => sig0000018f,
      I2 => start,
      I3 => sig00000198,
      I4 => NlwRenamedSig_OI_U0_i_synth_non_floating_point_arch_d_xfft_inst_FLOW_load_enable,
      O => sig00000184
    );
  blk0000100a : LUT3
    generic map(
      INIT => X"A8"
    )
    port map (
      I0 => ce,
      I1 => sig00000198,
      I2 => sig0000018f,
      O => sig00000185
    );
  blk0000100b : LUT4
    generic map(
      INIT => X"5504"
    )
    port map (
      I0 => sig00000187,
      I1 => sig0000018f,
      I2 => sig00000191,
      I3 => sig00000198,
      O => sig0000016e
    );
  blk0000100c : LUT2
    generic map(
      INIT => X"2"
    )
    port map (
      I0 => NlwRenamedSig_OI_xn_index(0),
      I1 => sig00000198,
      O => sig00000165
    );
  blk0000100d : LUT2
    generic map(
      INIT => X"2"
    )
    port map (
      I0 => NlwRenamedSig_OI_xn_index(1),
      I1 => sig00000198,
      O => sig00000164
    );
  blk0000100e : LUT2
    generic map(
      INIT => X"2"
    )
    port map (
      I0 => NlwRenamedSig_OI_xn_index(2),
      I1 => sig00000198,
      O => sig00000163
    );
  blk0000100f : LUT2
    generic map(
      INIT => X"2"
    )
    port map (
      I0 => NlwRenamedSig_OI_xn_index(3),
      I1 => sig00000198,
      O => sig00000162
    );
  blk00001010 : LUT2
    generic map(
      INIT => X"2"
    )
    port map (
      I0 => NlwRenamedSig_OI_xn_index(4),
      I1 => sig00000198,
      O => sig00000161
    );
  blk00001011 : LUT2
    generic map(
      INIT => X"4"
    )
    port map (
      I0 => sig00000198,
      I1 => NlwRenamedSig_OI_xn_index(5),
      O => sig00000160
    );
  blk00001012 : LUT2
    generic map(
      INIT => X"8"
    )
    port map (
      I0 => ce,
      I1 => sig00000190,
      O => sig00000168
    );
  blk00001013 : LUT2
    generic map(
      INIT => X"8"
    )
    port map (
      I0 => ce,
      I1 => cp_len_we,
      O => sig00000169
    );
  blk00001014 : LUT2
    generic map(
      INIT => X"8"
    )
    port map (
      I0 => ce,
      I1 => scale_sch_we,
      O => sig0000016a
    );
  blk00001015 : LUT2
    generic map(
      INIT => X"7"
    )
    port map (
      I0 => NlwRenamedSig_OI_rfs,
      I1 => start,
      O => sig0000016f
    );
  blk00001016 : LUT4
    generic map(
      INIT => X"F222"
    )
    port map (
      I0 => NlwRenamedSig_OI_U0_i_synth_non_floating_point_arch_d_xfft_inst_FLOW_load_enable,
      I1 => sig00000198,
      I2 => start,
      I3 => NlwRenamedSig_OI_rfs,
      O => sig00000170
    );
  blk00001017 : LUT3
    generic map(
      INIT => X"F8"
    )
    port map (
      I0 => sig00000189,
      I1 => sig0000018c,
      I2 => sig0000018d,
      O => sig00000176
    );
  blk00001018 : LUT2
    generic map(
      INIT => X"8"
    )
    port map (
      I0 => NlwRenamedSig_OI_U0_i_synth_non_floating_point_arch_d_xfft_inst_FLOW_load_enable,
      I1 => ce,
      O => sig00000186
    );
  blk00001019 : LUT4
    generic map(
      INIT => X"CC0A"
    )
    port map (
      I0 => sig00000192,
      I1 => sig0000011e,
      I2 => sig00000191,
      I3 => sig00000198,
      O => sig000001bf
    );
  blk0000101a : LUT4
    generic map(
      INIT => X"CC0A"
    )
    port map (
      I0 => sig00000193,
      I1 => sig0000011f,
      I2 => sig00000191,
      I3 => sig00000198,
      O => sig000001c0
    );
  blk0000101b : LUT4
    generic map(
      INIT => X"CC0A"
    )
    port map (
      I0 => sig00000194,
      I1 => sig00000120,
      I2 => sig00000191,
      I3 => sig00000198,
      O => sig000001c1
    );
  blk0000101c : LUT4
    generic map(
      INIT => X"CC0A"
    )
    port map (
      I0 => sig00000195,
      I1 => sig00000121,
      I2 => sig00000191,
      I3 => sig00000198,
      O => sig000001c2
    );
  blk0000101d : LUT4
    generic map(
      INIT => X"CC0A"
    )
    port map (
      I0 => sig00000196,
      I1 => sig00000122,
      I2 => sig00000191,
      I3 => sig00000198,
      O => sig000001c3
    );
  blk0000101e : LUT4
    generic map(
      INIT => X"BA10"
    )
    port map (
      I0 => sig00000198,
      I1 => sig00000191,
      I2 => sig00000197,
      I3 => sig00000123,
      O => sig000001c4
    );
  blk0000101f : LUT2
    generic map(
      INIT => X"B"
    )
    port map (
      I0 => sig00000198,
      I1 => sig00000191,
      O => sig000001be
    );
  blk00001020 : LUT4
    generic map(
      INIT => X"EA2A"
    )
    port map (
      I0 => sig0000025a,
      I1 => sig00000112,
      I2 => ce,
      I3 => sig0000011c,
      O => sig000001e9
    );
  blk00001021 : LUT3
    generic map(
      INIT => X"D8"
    )
    port map (
      I0 => ce,
      I1 => sig000001e7,
      I2 => sig000000ee,
      O => sig000001e8
    );
  blk00001022 : LUT2
    generic map(
      INIT => X"8"
    )
    port map (
      I0 => ce,
      I1 => sig00000282,
      O => sig000001ea
    );
  blk00001023 : LUT2
    generic map(
      INIT => X"2"
    )
    port map (
      I0 => sig00000283,
      I1 => sig000002a0,
      O => sig00000297
    );
  blk00001024 : LUT2
    generic map(
      INIT => X"2"
    )
    port map (
      I0 => sig00000284,
      I1 => sig000002a0,
      O => sig00000296
    );
  blk00001025 : LUT2
    generic map(
      INIT => X"2"
    )
    port map (
      I0 => sig00000285,
      I1 => sig000002a0,
      O => sig00000295
    );
  blk00001026 : LUT2
    generic map(
      INIT => X"4"
    )
    port map (
      I0 => sig000002a0,
      I1 => sig00000286,
      O => sig00000294
    );
  blk00001027 : LUT2
    generic map(
      INIT => X"4"
    )
    port map (
      I0 => sig000002a0,
      I1 => sig00000287,
      O => sig00000293
    );
  blk00001028 : LUT2
    generic map(
      INIT => X"4"
    )
    port map (
      I0 => sig000002a0,
      I1 => sig00000288,
      O => sig00000292
    );
  blk00001029 : LUT2
    generic map(
      INIT => X"8"
    )
    port map (
      I0 => sig0000029f,
      I1 => ce,
      O => sig0000029e
    );
  blk0000102a : LUT2
    generic map(
      INIT => X"2"
    )
    port map (
      I0 => sig0000027c,
      I1 => sig000002b8,
      O => sig000002af
    );
  blk0000102b : LUT2
    generic map(
      INIT => X"2"
    )
    port map (
      I0 => sig0000027d,
      I1 => sig000002b8,
      O => sig000002ae
    );
  blk0000102c : LUT2
    generic map(
      INIT => X"2"
    )
    port map (
      I0 => sig0000027e,
      I1 => sig000002b8,
      O => sig000002ad
    );
  blk0000102d : LUT2
    generic map(
      INIT => X"4"
    )
    port map (
      I0 => sig000002b8,
      I1 => sig0000027f,
      O => sig000002ac
    );
  blk0000102e : LUT2
    generic map(
      INIT => X"4"
    )
    port map (
      I0 => sig000002b8,
      I1 => sig00000280,
      O => sig000002ab
    );
  blk0000102f : LUT2
    generic map(
      INIT => X"4"
    )
    port map (
      I0 => sig000002b8,
      I1 => sig00000281,
      O => sig000002aa
    );
  blk00001030 : LUT2
    generic map(
      INIT => X"8"
    )
    port map (
      I0 => sig000002b7,
      I1 => ce,
      O => sig000002b6
    );
  blk00001031 : LUT4
    generic map(
      INIT => X"7D28"
    )
    port map (
      I0 => sig0000048e,
      I1 => sig0000026e,
      I2 => sig00000493,
      I3 => sig00000261,
      O => sig00000391
    );
  blk00001032 : LUT4
    generic map(
      INIT => X"7D28"
    )
    port map (
      I0 => sig0000048e,
      I1 => sig00000270,
      I2 => sig00000493,
      I3 => sig00000263,
      O => sig00000393
    );
  blk00001033 : LUT4
    generic map(
      INIT => X"7D28"
    )
    port map (
      I0 => sig0000048e,
      I1 => sig00000271,
      I2 => sig00000493,
      I3 => sig00000264,
      O => sig00000394
    );
  blk00001034 : LUT4
    generic map(
      INIT => X"7D28"
    )
    port map (
      I0 => sig0000048e,
      I1 => sig0000026f,
      I2 => sig00000493,
      I3 => sig00000262,
      O => sig00000392
    );
  blk00001035 : LUT4
    generic map(
      INIT => X"7D28"
    )
    port map (
      I0 => sig0000048e,
      I1 => sig00000272,
      I2 => sig00000493,
      I3 => sig00000265,
      O => sig00000395
    );
  blk00001036 : LUT4
    generic map(
      INIT => X"7D28"
    )
    port map (
      I0 => sig0000048e,
      I1 => sig00000273,
      I2 => sig00000493,
      I3 => sig00000266,
      O => sig00000396
    );
  blk00001037 : LUT4
    generic map(
      INIT => X"7D28"
    )
    port map (
      I0 => sig0000048e,
      I1 => sig00000275,
      I2 => sig00000493,
      I3 => sig00000268,
      O => sig00000398
    );
  blk00001038 : LUT4
    generic map(
      INIT => X"7D28"
    )
    port map (
      I0 => sig0000048e,
      I1 => sig00000276,
      I2 => sig00000493,
      I3 => sig00000269,
      O => sig00000399
    );
  blk00001039 : LUT4
    generic map(
      INIT => X"7D28"
    )
    port map (
      I0 => sig0000048e,
      I1 => sig00000274,
      I2 => sig00000493,
      I3 => sig00000267,
      O => sig00000397
    );
  blk0000103a : LUT4
    generic map(
      INIT => X"7D28"
    )
    port map (
      I0 => sig0000048e,
      I1 => sig00000278,
      I2 => sig00000493,
      I3 => sig0000026b,
      O => sig0000039b
    );
  blk0000103b : LUT4
    generic map(
      INIT => X"7D28"
    )
    port map (
      I0 => sig0000048e,
      I1 => sig00000279,
      I2 => sig00000493,
      I3 => sig0000026c,
      O => sig0000039c
    );
  blk0000103c : LUT4
    generic map(
      INIT => X"7D28"
    )
    port map (
      I0 => sig0000048e,
      I1 => sig00000277,
      I2 => sig00000493,
      I3 => sig0000026a,
      O => sig0000039a
    );
  blk0000103d : LUT4
    generic map(
      INIT => X"7D28"
    )
    port map (
      I0 => sig0000048e,
      I1 => sig0000027a,
      I2 => sig00000493,
      I3 => sig0000026d,
      O => sig0000039d
    );
  blk0000103e : LUT4
    generic map(
      INIT => X"D782"
    )
    port map (
      I0 => sig0000048e,
      I1 => sig00000261,
      I2 => sig00000493,
      I3 => sig0000026e,
      O => sig000003bb
    );
  blk0000103f : LUT4
    generic map(
      INIT => X"D782"
    )
    port map (
      I0 => sig0000048e,
      I1 => sig00000262,
      I2 => sig00000493,
      I3 => sig0000026f,
      O => sig000003bc
    );
  blk00001040 : LUT4
    generic map(
      INIT => X"D782"
    )
    port map (
      I0 => sig0000048e,
      I1 => sig00000263,
      I2 => sig00000493,
      I3 => sig00000270,
      O => sig000003bd
    );
  blk00001041 : LUT4
    generic map(
      INIT => X"D782"
    )
    port map (
      I0 => sig0000048e,
      I1 => sig00000265,
      I2 => sig00000493,
      I3 => sig00000272,
      O => sig000003bf
    );
  blk00001042 : LUT4
    generic map(
      INIT => X"D782"
    )
    port map (
      I0 => sig0000048e,
      I1 => sig00000266,
      I2 => sig00000493,
      I3 => sig00000273,
      O => sig000003c0
    );
  blk00001043 : LUT4
    generic map(
      INIT => X"D782"
    )
    port map (
      I0 => sig0000048e,
      I1 => sig00000264,
      I2 => sig00000493,
      I3 => sig00000271,
      O => sig000003be
    );
  blk00001044 : LUT4
    generic map(
      INIT => X"D782"
    )
    port map (
      I0 => sig0000048e,
      I1 => sig00000268,
      I2 => sig00000493,
      I3 => sig00000275,
      O => sig000003c2
    );
  blk00001045 : LUT4
    generic map(
      INIT => X"D782"
    )
    port map (
      I0 => sig0000048e,
      I1 => sig00000269,
      I2 => sig00000493,
      I3 => sig00000276,
      O => sig000003c3
    );
  blk00001046 : LUT4
    generic map(
      INIT => X"D782"
    )
    port map (
      I0 => sig0000048e,
      I1 => sig00000267,
      I2 => sig00000493,
      I3 => sig00000274,
      O => sig000003c1
    );
  blk00001047 : LUT4
    generic map(
      INIT => X"D782"
    )
    port map (
      I0 => sig0000048e,
      I1 => sig0000026b,
      I2 => sig00000493,
      I3 => sig00000278,
      O => sig000003c5
    );
  blk00001048 : LUT4
    generic map(
      INIT => X"D782"
    )
    port map (
      I0 => sig0000048e,
      I1 => sig0000026c,
      I2 => sig00000493,
      I3 => sig00000279,
      O => sig000003c6
    );
  blk00001049 : LUT4
    generic map(
      INIT => X"D782"
    )
    port map (
      I0 => sig0000048e,
      I1 => sig0000026a,
      I2 => sig00000493,
      I3 => sig00000277,
      O => sig000003c4
    );
  blk0000104a : LUT4
    generic map(
      INIT => X"D782"
    )
    port map (
      I0 => sig0000048e,
      I1 => sig0000026d,
      I2 => sig00000493,
      I3 => sig0000027a,
      O => sig000003c7
    );
  blk0000104b : LUT3
    generic map(
      INIT => X"D8"
    )
    port map (
      I0 => sig0000048f,
      I1 => sig0000041c,
      I2 => sig00000438,
      O => sig00000376
    );
  blk0000104c : LUT3
    generic map(
      INIT => X"D8"
    )
    port map (
      I0 => sig0000048f,
      I1 => sig0000041b,
      I2 => sig00000437,
      O => sig00000377
    );
  blk0000104d : LUT3
    generic map(
      INIT => X"D8"
    )
    port map (
      I0 => sig0000048f,
      I1 => sig0000041d,
      I2 => sig00000439,
      O => sig00000375
    );
  blk0000104e : LUT3
    generic map(
      INIT => X"D8"
    )
    port map (
      I0 => sig0000048f,
      I1 => sig0000041a,
      I2 => sig00000436,
      O => sig00000378
    );
  blk0000104f : LUT3
    generic map(
      INIT => X"D8"
    )
    port map (
      I0 => sig0000048f,
      I1 => sig00000419,
      I2 => sig00000435,
      O => sig00000379
    );
  blk00001050 : LUT3
    generic map(
      INIT => X"D8"
    )
    port map (
      I0 => sig0000048f,
      I1 => sig00000417,
      I2 => sig00000433,
      O => sig0000037b
    );
  blk00001051 : LUT3
    generic map(
      INIT => X"D8"
    )
    port map (
      I0 => sig0000048f,
      I1 => sig00000416,
      I2 => sig00000432,
      O => sig0000037c
    );
  blk00001052 : LUT3
    generic map(
      INIT => X"D8"
    )
    port map (
      I0 => sig0000048f,
      I1 => sig00000418,
      I2 => sig00000434,
      O => sig0000037a
    );
  blk00001053 : LUT3
    generic map(
      INIT => X"D8"
    )
    port map (
      I0 => sig0000048f,
      I1 => sig00000414,
      I2 => sig00000430,
      O => sig0000037e
    );
  blk00001054 : LUT3
    generic map(
      INIT => X"D8"
    )
    port map (
      I0 => sig0000048f,
      I1 => sig00000413,
      I2 => sig0000042f,
      O => sig0000037f
    );
  blk00001055 : LUT3
    generic map(
      INIT => X"D8"
    )
    port map (
      I0 => sig0000048f,
      I1 => sig00000415,
      I2 => sig00000431,
      O => sig0000037d
    );
  blk00001056 : LUT3
    generic map(
      INIT => X"D8"
    )
    port map (
      I0 => sig0000048f,
      I1 => sig00000411,
      I2 => sig0000042d,
      O => sig00000381
    );
  blk00001057 : LUT3
    generic map(
      INIT => X"D8"
    )
    port map (
      I0 => sig0000048f,
      I1 => sig00000410,
      I2 => sig0000042c,
      O => sig00000382
    );
  blk00001058 : LUT3
    generic map(
      INIT => X"D8"
    )
    port map (
      I0 => sig0000048f,
      I1 => sig00000412,
      I2 => sig0000042e,
      O => sig00000380
    );
  blk00001059 : LUT3
    generic map(
      INIT => X"D8"
    )
    port map (
      I0 => sig0000048f,
      I1 => sig00000439,
      I2 => sig0000041d,
      O => sig00000383
    );
  blk0000105a : LUT3
    generic map(
      INIT => X"D8"
    )
    port map (
      I0 => sig0000048f,
      I1 => sig00000438,
      I2 => sig0000041c,
      O => sig00000384
    );
  blk0000105b : LUT3
    generic map(
      INIT => X"D8"
    )
    port map (
      I0 => sig0000048f,
      I1 => sig00000436,
      I2 => sig0000041a,
      O => sig00000386
    );
  blk0000105c : LUT3
    generic map(
      INIT => X"D8"
    )
    port map (
      I0 => sig0000048f,
      I1 => sig00000435,
      I2 => sig00000419,
      O => sig00000387
    );
  blk0000105d : LUT3
    generic map(
      INIT => X"D8"
    )
    port map (
      I0 => sig0000048f,
      I1 => sig00000437,
      I2 => sig0000041b,
      O => sig00000385
    );
  blk0000105e : LUT3
    generic map(
      INIT => X"D8"
    )
    port map (
      I0 => sig0000048f,
      I1 => sig00000433,
      I2 => sig00000417,
      O => sig00000389
    );
  blk0000105f : LUT3
    generic map(
      INIT => X"D8"
    )
    port map (
      I0 => sig0000048f,
      I1 => sig00000432,
      I2 => sig00000416,
      O => sig0000038a
    );
  blk00001060 : LUT3
    generic map(
      INIT => X"D8"
    )
    port map (
      I0 => sig0000048f,
      I1 => sig00000434,
      I2 => sig00000418,
      O => sig00000388
    );
  blk00001061 : LUT3
    generic map(
      INIT => X"D8"
    )
    port map (
      I0 => sig0000048f,
      I1 => sig00000430,
      I2 => sig00000414,
      O => sig0000038c
    );
  blk00001062 : LUT3
    generic map(
      INIT => X"D8"
    )
    port map (
      I0 => sig0000048f,
      I1 => sig0000042f,
      I2 => sig00000413,
      O => sig0000038d
    );
  blk00001063 : LUT3
    generic map(
      INIT => X"D8"
    )
    port map (
      I0 => sig0000048f,
      I1 => sig00000431,
      I2 => sig00000415,
      O => sig0000038b
    );
  blk00001064 : LUT3
    generic map(
      INIT => X"D8"
    )
    port map (
      I0 => sig0000048f,
      I1 => sig0000042e,
      I2 => sig00000412,
      O => sig0000038e
    );
  blk00001065 : LUT3
    generic map(
      INIT => X"D8"
    )
    port map (
      I0 => sig0000048f,
      I1 => sig0000042d,
      I2 => sig00000411,
      O => sig0000038f
    );
  blk00001066 : LUT3
    generic map(
      INIT => X"D8"
    )
    port map (
      I0 => sig0000048f,
      I1 => sig0000042c,
      I2 => sig00000410,
      O => sig00000390
    );
  blk00001067 : LUT3
    generic map(
      INIT => X"D8"
    )
    port map (
      I0 => sig00000491,
      I1 => sig00000462,
      I2 => sig000003f2,
      O => sig0000035a
    );
  blk00001068 : LUT3
    generic map(
      INIT => X"D8"
    )
    port map (
      I0 => sig00000491,
      I1 => sig00000461,
      I2 => sig000003f1,
      O => sig0000035b
    );
  blk00001069 : LUT3
    generic map(
      INIT => X"D8"
    )
    port map (
      I0 => sig00000491,
      I1 => sig00000463,
      I2 => sig000003f3,
      O => sig00000359
    );
  blk0000106a : LUT3
    generic map(
      INIT => X"D8"
    )
    port map (
      I0 => sig00000491,
      I1 => sig0000045f,
      I2 => sig000003ef,
      O => sig0000035d
    );
  blk0000106b : LUT3
    generic map(
      INIT => X"D8"
    )
    port map (
      I0 => sig00000491,
      I1 => sig0000045e,
      I2 => sig000003ee,
      O => sig0000035e
    );
  blk0000106c : LUT3
    generic map(
      INIT => X"D8"
    )
    port map (
      I0 => sig00000491,
      I1 => sig00000460,
      I2 => sig000003f0,
      O => sig0000035c
    );
  blk0000106d : LUT3
    generic map(
      INIT => X"D8"
    )
    port map (
      I0 => sig00000491,
      I1 => sig0000045c,
      I2 => sig000003ec,
      O => sig00000360
    );
  blk0000106e : LUT3
    generic map(
      INIT => X"D8"
    )
    port map (
      I0 => sig00000491,
      I1 => sig0000045b,
      I2 => sig000003eb,
      O => sig00000361
    );
  blk0000106f : LUT3
    generic map(
      INIT => X"D8"
    )
    port map (
      I0 => sig00000491,
      I1 => sig0000045d,
      I2 => sig000003ed,
      O => sig0000035f
    );
  blk00001070 : LUT3
    generic map(
      INIT => X"D8"
    )
    port map (
      I0 => sig00000491,
      I1 => sig0000045a,
      I2 => sig000003ea,
      O => sig00000362
    );
  blk00001071 : LUT3
    generic map(
      INIT => X"D8"
    )
    port map (
      I0 => sig00000491,
      I1 => sig00000459,
      I2 => sig000003e9,
      O => sig00000363
    );
  blk00001072 : LUT3
    generic map(
      INIT => X"D8"
    )
    port map (
      I0 => sig00000491,
      I1 => sig00000457,
      I2 => sig000003e7,
      O => sig00000365
    );
  blk00001073 : LUT3
    generic map(
      INIT => X"D8"
    )
    port map (
      I0 => sig00000491,
      I1 => sig00000456,
      I2 => sig000003e6,
      O => sig00000366
    );
  blk00001074 : LUT3
    generic map(
      INIT => X"D8"
    )
    port map (
      I0 => sig00000491,
      I1 => sig00000458,
      I2 => sig000003e8,
      O => sig00000364
    );
  blk00001075 : LUT3
    generic map(
      INIT => X"D8"
    )
    port map (
      I0 => sig00000491,
      I1 => sig000003f2,
      I2 => sig00000462,
      O => sig00000368
    );
  blk00001076 : LUT3
    generic map(
      INIT => X"D8"
    )
    port map (
      I0 => sig00000491,
      I1 => sig000003f1,
      I2 => sig00000461,
      O => sig00000369
    );
  blk00001077 : LUT3
    generic map(
      INIT => X"D8"
    )
    port map (
      I0 => sig00000491,
      I1 => sig000003f3,
      I2 => sig00000463,
      O => sig00000367
    );
  blk00001078 : LUT3
    generic map(
      INIT => X"D8"
    )
    port map (
      I0 => sig00000491,
      I1 => sig000003ef,
      I2 => sig0000045f,
      O => sig0000036b
    );
  blk00001079 : LUT3
    generic map(
      INIT => X"D8"
    )
    port map (
      I0 => sig00000491,
      I1 => sig000003ee,
      I2 => sig0000045e,
      O => sig0000036c
    );
  blk0000107a : LUT3
    generic map(
      INIT => X"D8"
    )
    port map (
      I0 => sig00000491,
      I1 => sig000003f0,
      I2 => sig00000460,
      O => sig0000036a
    );
  blk0000107b : LUT3
    generic map(
      INIT => X"D8"
    )
    port map (
      I0 => sig00000491,
      I1 => sig000003ed,
      I2 => sig0000045d,
      O => sig0000036d
    );
  blk0000107c : LUT3
    generic map(
      INIT => X"D8"
    )
    port map (
      I0 => sig00000491,
      I1 => sig000003ec,
      I2 => sig0000045c,
      O => sig0000036e
    );
  blk0000107d : LUT3
    generic map(
      INIT => X"D8"
    )
    port map (
      I0 => sig00000491,
      I1 => sig000003ea,
      I2 => sig0000045a,
      O => sig00000370
    );
  blk0000107e : LUT3
    generic map(
      INIT => X"D8"
    )
    port map (
      I0 => sig00000491,
      I1 => sig000003e9,
      I2 => sig00000459,
      O => sig00000371
    );
  blk0000107f : LUT3
    generic map(
      INIT => X"D8"
    )
    port map (
      I0 => sig00000491,
      I1 => sig000003eb,
      I2 => sig0000045b,
      O => sig0000036f
    );
  blk00001080 : LUT3
    generic map(
      INIT => X"D8"
    )
    port map (
      I0 => sig00000491,
      I1 => sig000003e7,
      I2 => sig00000457,
      O => sig00000373
    );
  blk00001081 : LUT3
    generic map(
      INIT => X"D8"
    )
    port map (
      I0 => sig00000491,
      I1 => sig000003e6,
      I2 => sig00000456,
      O => sig00000374
    );
  blk00001082 : LUT3
    generic map(
      INIT => X"D8"
    )
    port map (
      I0 => sig00000491,
      I1 => sig000003e8,
      I2 => sig00000458,
      O => sig00000372
    );
  blk00001083 : LUT2
    generic map(
      INIT => X"8"
    )
    port map (
      I0 => sig0000048e,
      I1 => sig00000493,
      O => sig0000039e
    );
  blk00001084 : LUT2
    generic map(
      INIT => X"4"
    )
    port map (
      I0 => sig00000493,
      I1 => sig0000048e,
      O => sig000003c8
    );
  blk00001085 : LUT2
    generic map(
      INIT => X"8"
    )
    port map (
      I0 => sig00000250,
      I1 => sig0000024f,
      O => sig000003e5
    );
  blk00001086 : LUT4
    generic map(
      INIT => X"EA2A"
    )
    port map (
      I0 => sig00000a60,
      I1 => sig000000ee,
      I2 => ce,
      I3 => sig000000ed,
      O => sig000009f7
    );
  blk00001087 : LUT3
    generic map(
      INIT => X"D8"
    )
    port map (
      I0 => ce,
      I1 => sig000009f5,
      I2 => sig000000ca,
      O => sig000009f6
    );
  blk00001088 : LUT2
    generic map(
      INIT => X"8"
    )
    port map (
      I0 => ce,
      I1 => sig00000a86,
      O => sig000009f8
    );
  blk00001089 : LUT2
    generic map(
      INIT => X"2"
    )
    port map (
      I0 => sig00000a87,
      I1 => sig00000aa2,
      O => sig00000a99
    );
  blk0000108a : LUT2
    generic map(
      INIT => X"2"
    )
    port map (
      I0 => sig00000a88,
      I1 => sig00000aa2,
      O => sig00000a98
    );
  blk0000108b : LUT2
    generic map(
      INIT => X"2"
    )
    port map (
      I0 => sig00000a89,
      I1 => sig00000aa2,
      O => sig00000a97
    );
  blk0000108c : LUT2
    generic map(
      INIT => X"4"
    )
    port map (
      I0 => sig00000aa2,
      I1 => sig00000a8a,
      O => sig00000a96
    );
  blk0000108d : LUT2
    generic map(
      INIT => X"4"
    )
    port map (
      I0 => sig00000aa2,
      I1 => sig00000aa3,
      O => sig00000a95
    );
  blk0000108e : LUT2
    generic map(
      INIT => X"4"
    )
    port map (
      I0 => sig00000aa2,
      I1 => sig00000aa4,
      O => sig00000a94
    );
  blk0000108f : LUT2
    generic map(
      INIT => X"8"
    )
    port map (
      I0 => sig00000aa1,
      I1 => ce,
      O => sig00000aa0
    );
  blk00001090 : LUT2
    generic map(
      INIT => X"4"
    )
    port map (
      I0 => sig00000abc,
      I1 => sig00000a82,
      O => sig00000ab3
    );
  blk00001091 : LUT2
    generic map(
      INIT => X"4"
    )
    port map (
      I0 => sig00000abc,
      I1 => sig00000a83,
      O => sig00000ab2
    );
  blk00001092 : LUT2
    generic map(
      INIT => X"2"
    )
    port map (
      I0 => sig00000a84,
      I1 => sig00000abc,
      O => sig00000ab1
    );
  blk00001093 : LUT2
    generic map(
      INIT => X"4"
    )
    port map (
      I0 => sig00000abc,
      I1 => sig00000a85,
      O => sig00000ab0
    );
  blk00001094 : LUT2
    generic map(
      INIT => X"4"
    )
    port map (
      I0 => sig00000abc,
      I1 => sig00000abd,
      O => sig00000aaf
    );
  blk00001095 : LUT2
    generic map(
      INIT => X"4"
    )
    port map (
      I0 => sig00000abc,
      I1 => sig00000abe,
      O => sig00000aae
    );
  blk00001096 : LUT2
    generic map(
      INIT => X"8"
    )
    port map (
      I0 => sig00000abb,
      I1 => ce,
      O => sig00000aba
    );
  blk00001097 : LUT3
    generic map(
      INIT => X"D8"
    )
    port map (
      I0 => sig00000b31,
      I1 => sig00000b09,
      I2 => sig00000b23,
      O => sig00000ac0
    );
  blk00001098 : LUT3
    generic map(
      INIT => X"D8"
    )
    port map (
      I0 => sig00000b31,
      I1 => sig00000b08,
      I2 => sig00000b22,
      O => sig00000ac1
    );
  blk00001099 : LUT3
    generic map(
      INIT => X"D8"
    )
    port map (
      I0 => sig00000b31,
      I1 => sig00000b0a,
      I2 => sig00000b24,
      O => sig00000abf
    );
  blk0000109a : LUT3
    generic map(
      INIT => X"D8"
    )
    port map (
      I0 => sig00000b31,
      I1 => sig00000b07,
      I2 => sig00000b21,
      O => sig00000ac2
    );
  blk0000109b : LUT3
    generic map(
      INIT => X"D8"
    )
    port map (
      I0 => sig00000b31,
      I1 => sig00000b06,
      I2 => sig00000b20,
      O => sig00000ac3
    );
  blk0000109c : LUT3
    generic map(
      INIT => X"D8"
    )
    port map (
      I0 => sig00000b31,
      I1 => sig00000b05,
      I2 => sig00000b1f,
      O => sig00000ac4
    );
  blk0000109d : LUT3
    generic map(
      INIT => X"D8"
    )
    port map (
      I0 => sig00000b31,
      I1 => sig00000b04,
      I2 => sig00000b1e,
      O => sig00000ac5
    );
  blk0000109e : LUT3
    generic map(
      INIT => X"D8"
    )
    port map (
      I0 => sig00000b31,
      I1 => sig00000b02,
      I2 => sig00000b1c,
      O => sig00000ac7
    );
  blk0000109f : LUT3
    generic map(
      INIT => X"D8"
    )
    port map (
      I0 => sig00000b31,
      I1 => sig00000b01,
      I2 => sig00000b1b,
      O => sig00000ac8
    );
  blk000010a0 : LUT3
    generic map(
      INIT => X"D8"
    )
    port map (
      I0 => sig00000b31,
      I1 => sig00000b03,
      I2 => sig00000b1d,
      O => sig00000ac6
    );
  blk000010a1 : LUT3
    generic map(
      INIT => X"D8"
    )
    port map (
      I0 => sig00000b31,
      I1 => sig00000b00,
      I2 => sig00000b1a,
      O => sig00000ac9
    );
  blk000010a2 : LUT3
    generic map(
      INIT => X"D8"
    )
    port map (
      I0 => sig00000b31,
      I1 => sig00000aff,
      I2 => sig00000b19,
      O => sig00000aca
    );
  blk000010a3 : LUT3
    generic map(
      INIT => X"D8"
    )
    port map (
      I0 => sig00000b31,
      I1 => sig00000afe,
      I2 => sig00000b18,
      O => sig00000acb
    );
  blk000010a4 : LUT3
    generic map(
      INIT => X"D8"
    )
    port map (
      I0 => sig00000b31,
      I1 => sig00000b24,
      I2 => sig00000b0a,
      O => sig00000acc
    );
  blk000010a5 : LUT3
    generic map(
      INIT => X"D8"
    )
    port map (
      I0 => sig00000b31,
      I1 => sig00000b22,
      I2 => sig00000b08,
      O => sig00000ace
    );
  blk000010a6 : LUT3
    generic map(
      INIT => X"D8"
    )
    port map (
      I0 => sig00000b31,
      I1 => sig00000b21,
      I2 => sig00000b07,
      O => sig00000acf
    );
  blk000010a7 : LUT3
    generic map(
      INIT => X"D8"
    )
    port map (
      I0 => sig00000b31,
      I1 => sig00000b23,
      I2 => sig00000b09,
      O => sig00000acd
    );
  blk000010a8 : LUT3
    generic map(
      INIT => X"D8"
    )
    port map (
      I0 => sig00000b31,
      I1 => sig00000b20,
      I2 => sig00000b06,
      O => sig00000ad0
    );
  blk000010a9 : LUT3
    generic map(
      INIT => X"D8"
    )
    port map (
      I0 => sig00000b31,
      I1 => sig00000b1f,
      I2 => sig00000b05,
      O => sig00000ad1
    );
  blk000010aa : LUT3
    generic map(
      INIT => X"D8"
    )
    port map (
      I0 => sig00000b31,
      I1 => sig00000b1e,
      I2 => sig00000b04,
      O => sig00000ad2
    );
  blk000010ab : LUT3
    generic map(
      INIT => X"D8"
    )
    port map (
      I0 => sig00000b31,
      I1 => sig00000b1d,
      I2 => sig00000b03,
      O => sig00000ad3
    );
  blk000010ac : LUT3
    generic map(
      INIT => X"D8"
    )
    port map (
      I0 => sig00000b31,
      I1 => sig00000b1b,
      I2 => sig00000b01,
      O => sig00000ad5
    );
  blk000010ad : LUT3
    generic map(
      INIT => X"D8"
    )
    port map (
      I0 => sig00000b31,
      I1 => sig00000b1a,
      I2 => sig00000b00,
      O => sig00000ad6
    );
  blk000010ae : LUT3
    generic map(
      INIT => X"D8"
    )
    port map (
      I0 => sig00000b31,
      I1 => sig00000b1c,
      I2 => sig00000b02,
      O => sig00000ad4
    );
  blk000010af : LUT3
    generic map(
      INIT => X"D8"
    )
    port map (
      I0 => sig00000b31,
      I1 => sig00000b19,
      I2 => sig00000aff,
      O => sig00000ad7
    );
  blk000010b0 : LUT3
    generic map(
      INIT => X"D8"
    )
    port map (
      I0 => sig00000b31,
      I1 => sig00000b18,
      I2 => sig00000afe,
      O => sig00000ad8
    );
  blk000010b1 : LUT3
    generic map(
      INIT => X"D8"
    )
    port map (
      I0 => sig00000111,
      I1 => sig00000b3f,
      I2 => sig00000106,
      O => sig00000ad9
    );
  blk000010b2 : LUT3
    generic map(
      INIT => X"D8"
    )
    port map (
      I0 => sig00000111,
      I1 => sig00000b3e,
      I2 => sig00000105,
      O => sig00000ada
    );
  blk000010b3 : LUT3
    generic map(
      INIT => X"D8"
    )
    port map (
      I0 => sig00000111,
      I1 => sig00000b3c,
      I2 => sig00000103,
      O => sig00000adc
    );
  blk000010b4 : LUT3
    generic map(
      INIT => X"D8"
    )
    port map (
      I0 => sig00000111,
      I1 => sig00000b3b,
      I2 => sig00000102,
      O => sig00000add
    );
  blk000010b5 : LUT3
    generic map(
      INIT => X"D8"
    )
    port map (
      I0 => sig00000111,
      I1 => sig00000b3d,
      I2 => sig00000104,
      O => sig00000adb
    );
  blk000010b6 : LUT3
    generic map(
      INIT => X"D8"
    )
    port map (
      I0 => sig00000111,
      I1 => sig00000b3a,
      I2 => sig00000101,
      O => sig00000ade
    );
  blk000010b7 : LUT3
    generic map(
      INIT => X"D8"
    )
    port map (
      I0 => sig00000111,
      I1 => sig00000b39,
      I2 => sig00000100,
      O => sig00000adf
    );
  blk000010b8 : LUT3
    generic map(
      INIT => X"D8"
    )
    port map (
      I0 => sig00000111,
      I1 => sig00000b38,
      I2 => sig000000ff,
      O => sig00000ae0
    );
  blk000010b9 : LUT3
    generic map(
      INIT => X"D8"
    )
    port map (
      I0 => sig00000111,
      I1 => sig00000b37,
      I2 => sig000000fe,
      O => sig00000ae1
    );
  blk000010ba : LUT3
    generic map(
      INIT => X"D8"
    )
    port map (
      I0 => sig00000111,
      I1 => sig00000b35,
      I2 => sig000000fc,
      O => sig00000ae3
    );
  blk000010bb : LUT3
    generic map(
      INIT => X"D8"
    )
    port map (
      I0 => sig00000111,
      I1 => sig00000b34,
      I2 => sig000000fb,
      O => sig00000ae4
    );
  blk000010bc : LUT3
    generic map(
      INIT => X"D8"
    )
    port map (
      I0 => sig00000111,
      I1 => sig00000b36,
      I2 => sig000000fd,
      O => sig00000ae2
    );
  blk000010bd : LUT3
    generic map(
      INIT => X"D8"
    )
    port map (
      I0 => sig00000111,
      I1 => sig00000106,
      I2 => sig00000b3f,
      O => sig00000ae5
    );
  blk000010be : LUT3
    generic map(
      INIT => X"D8"
    )
    port map (
      I0 => sig00000111,
      I1 => sig00000105,
      I2 => sig00000b3e,
      O => sig00000ae6
    );
  blk000010bf : LUT3
    generic map(
      INIT => X"D8"
    )
    port map (
      I0 => sig00000111,
      I1 => sig00000104,
      I2 => sig00000b3d,
      O => sig00000ae7
    );
  blk000010c0 : LUT3
    generic map(
      INIT => X"D8"
    )
    port map (
      I0 => sig00000111,
      I1 => sig00000103,
      I2 => sig00000b3c,
      O => sig00000ae8
    );
  blk000010c1 : LUT3
    generic map(
      INIT => X"D8"
    )
    port map (
      I0 => sig00000111,
      I1 => sig00000102,
      I2 => sig00000b3b,
      O => sig00000ae9
    );
  blk000010c2 : LUT3
    generic map(
      INIT => X"D8"
    )
    port map (
      I0 => sig00000111,
      I1 => sig00000101,
      I2 => sig00000b3a,
      O => sig00000aea
    );
  blk000010c3 : LUT3
    generic map(
      INIT => X"D8"
    )
    port map (
      I0 => sig00000111,
      I1 => sig00000100,
      I2 => sig00000b39,
      O => sig00000aeb
    );
  blk000010c4 : LUT3
    generic map(
      INIT => X"D8"
    )
    port map (
      I0 => sig00000111,
      I1 => sig000000ff,
      I2 => sig00000b38,
      O => sig00000aec
    );
  blk000010c5 : LUT3
    generic map(
      INIT => X"D8"
    )
    port map (
      I0 => sig00000111,
      I1 => sig000000fe,
      I2 => sig00000b37,
      O => sig00000aed
    );
  blk000010c6 : LUT3
    generic map(
      INIT => X"D8"
    )
    port map (
      I0 => sig00000111,
      I1 => sig000000fd,
      I2 => sig00000b36,
      O => sig00000aee
    );
  blk000010c7 : LUT3
    generic map(
      INIT => X"D8"
    )
    port map (
      I0 => sig00000111,
      I1 => sig000000fc,
      I2 => sig00000b35,
      O => sig00000aef
    );
  blk000010c8 : LUT3
    generic map(
      INIT => X"D8"
    )
    port map (
      I0 => sig00000111,
      I1 => sig000000fb,
      I2 => sig00000b34,
      O => sig00000af0
    );
  blk000010c9 : LUT4
    generic map(
      INIT => X"7D28"
    )
    port map (
      I0 => sig00000c8d,
      I1 => sig00000a74,
      I2 => sig00000c92,
      I3 => sig00000a67,
      O => sig00000b90
    );
  blk000010ca : LUT4
    generic map(
      INIT => X"7D28"
    )
    port map (
      I0 => sig00000c8d,
      I1 => sig00000a76,
      I2 => sig00000c92,
      I3 => sig00000a69,
      O => sig00000b92
    );
  blk000010cb : LUT4
    generic map(
      INIT => X"7D28"
    )
    port map (
      I0 => sig00000c8d,
      I1 => sig00000a77,
      I2 => sig00000c92,
      I3 => sig00000a6a,
      O => sig00000b93
    );
  blk000010cc : LUT4
    generic map(
      INIT => X"7D28"
    )
    port map (
      I0 => sig00000c8d,
      I1 => sig00000a75,
      I2 => sig00000c92,
      I3 => sig00000a68,
      O => sig00000b91
    );
  blk000010cd : LUT4
    generic map(
      INIT => X"7D28"
    )
    port map (
      I0 => sig00000c8d,
      I1 => sig00000a78,
      I2 => sig00000c92,
      I3 => sig00000a6b,
      O => sig00000b94
    );
  blk000010ce : LUT4
    generic map(
      INIT => X"7D28"
    )
    port map (
      I0 => sig00000c8d,
      I1 => sig00000a79,
      I2 => sig00000c92,
      I3 => sig00000a6c,
      O => sig00000b95
    );
  blk000010cf : LUT4
    generic map(
      INIT => X"7D28"
    )
    port map (
      I0 => sig00000c8d,
      I1 => sig00000a7b,
      I2 => sig00000c92,
      I3 => sig00000a6e,
      O => sig00000b97
    );
  blk000010d0 : LUT4
    generic map(
      INIT => X"7D28"
    )
    port map (
      I0 => sig00000c8d,
      I1 => sig00000a7c,
      I2 => sig00000c92,
      I3 => sig00000a6f,
      O => sig00000b98
    );
  blk000010d1 : LUT4
    generic map(
      INIT => X"7D28"
    )
    port map (
      I0 => sig00000c8d,
      I1 => sig00000a7a,
      I2 => sig00000c92,
      I3 => sig00000a6d,
      O => sig00000b96
    );
  blk000010d2 : LUT4
    generic map(
      INIT => X"7D28"
    )
    port map (
      I0 => sig00000c8d,
      I1 => sig00000a7e,
      I2 => sig00000c92,
      I3 => sig00000a71,
      O => sig00000b9a
    );
  blk000010d3 : LUT4
    generic map(
      INIT => X"7D28"
    )
    port map (
      I0 => sig00000c8d,
      I1 => sig00000a7f,
      I2 => sig00000c92,
      I3 => sig00000a72,
      O => sig00000b9b
    );
  blk000010d4 : LUT4
    generic map(
      INIT => X"7D28"
    )
    port map (
      I0 => sig00000c8d,
      I1 => sig00000a7d,
      I2 => sig00000c92,
      I3 => sig00000a70,
      O => sig00000b99
    );
  blk000010d5 : LUT4
    generic map(
      INIT => X"7D28"
    )
    port map (
      I0 => sig00000c8d,
      I1 => sig00000a80,
      I2 => sig00000c92,
      I3 => sig00000a73,
      O => sig00000b9c
    );
  blk000010d6 : LUT4
    generic map(
      INIT => X"D782"
    )
    port map (
      I0 => sig00000c8d,
      I1 => sig00000a67,
      I2 => sig00000c92,
      I3 => sig00000a74,
      O => sig00000bba
    );
  blk000010d7 : LUT4
    generic map(
      INIT => X"D782"
    )
    port map (
      I0 => sig00000c8d,
      I1 => sig00000a68,
      I2 => sig00000c92,
      I3 => sig00000a75,
      O => sig00000bbb
    );
  blk000010d8 : LUT4
    generic map(
      INIT => X"D782"
    )
    port map (
      I0 => sig00000c8d,
      I1 => sig00000a69,
      I2 => sig00000c92,
      I3 => sig00000a76,
      O => sig00000bbc
    );
  blk000010d9 : LUT4
    generic map(
      INIT => X"D782"
    )
    port map (
      I0 => sig00000c8d,
      I1 => sig00000a6b,
      I2 => sig00000c92,
      I3 => sig00000a78,
      O => sig00000bbe
    );
  blk000010da : LUT4
    generic map(
      INIT => X"D782"
    )
    port map (
      I0 => sig00000c8d,
      I1 => sig00000a6c,
      I2 => sig00000c92,
      I3 => sig00000a79,
      O => sig00000bbf
    );
  blk000010db : LUT4
    generic map(
      INIT => X"D782"
    )
    port map (
      I0 => sig00000c8d,
      I1 => sig00000a6a,
      I2 => sig00000c92,
      I3 => sig00000a77,
      O => sig00000bbd
    );
  blk000010dc : LUT4
    generic map(
      INIT => X"D782"
    )
    port map (
      I0 => sig00000c8d,
      I1 => sig00000a6e,
      I2 => sig00000c92,
      I3 => sig00000a7b,
      O => sig00000bc1
    );
  blk000010dd : LUT4
    generic map(
      INIT => X"D782"
    )
    port map (
      I0 => sig00000c8d,
      I1 => sig00000a6f,
      I2 => sig00000c92,
      I3 => sig00000a7c,
      O => sig00000bc2
    );
  blk000010de : LUT4
    generic map(
      INIT => X"D782"
    )
    port map (
      I0 => sig00000c8d,
      I1 => sig00000a6d,
      I2 => sig00000c92,
      I3 => sig00000a7a,
      O => sig00000bc0
    );
  blk000010df : LUT4
    generic map(
      INIT => X"D782"
    )
    port map (
      I0 => sig00000c8d,
      I1 => sig00000a71,
      I2 => sig00000c92,
      I3 => sig00000a7e,
      O => sig00000bc4
    );
  blk000010e0 : LUT4
    generic map(
      INIT => X"D782"
    )
    port map (
      I0 => sig00000c8d,
      I1 => sig00000a72,
      I2 => sig00000c92,
      I3 => sig00000a7f,
      O => sig00000bc5
    );
  blk000010e1 : LUT4
    generic map(
      INIT => X"D782"
    )
    port map (
      I0 => sig00000c8d,
      I1 => sig00000a70,
      I2 => sig00000c92,
      I3 => sig00000a7d,
      O => sig00000bc3
    );
  blk000010e2 : LUT4
    generic map(
      INIT => X"D782"
    )
    port map (
      I0 => sig00000c8d,
      I1 => sig00000a73,
      I2 => sig00000c92,
      I3 => sig00000a80,
      O => sig00000bc6
    );
  blk000010e3 : LUT3
    generic map(
      INIT => X"D8"
    )
    port map (
      I0 => sig00000c8e,
      I1 => sig00000c1c,
      I2 => sig00000c38,
      O => sig00000b74
    );
  blk000010e4 : LUT3
    generic map(
      INIT => X"D8"
    )
    port map (
      I0 => sig00000c8e,
      I1 => sig00000c1a,
      I2 => sig00000c36,
      O => sig00000b76
    );
  blk000010e5 : LUT3
    generic map(
      INIT => X"D8"
    )
    port map (
      I0 => sig00000c8e,
      I1 => sig00000c19,
      I2 => sig00000c35,
      O => sig00000b77
    );
  blk000010e6 : LUT3
    generic map(
      INIT => X"D8"
    )
    port map (
      I0 => sig00000c8e,
      I1 => sig00000c1b,
      I2 => sig00000c37,
      O => sig00000b75
    );
  blk000010e7 : LUT3
    generic map(
      INIT => X"D8"
    )
    port map (
      I0 => sig00000c8e,
      I1 => sig00000c17,
      I2 => sig00000c33,
      O => sig00000b79
    );
  blk000010e8 : LUT3
    generic map(
      INIT => X"D8"
    )
    port map (
      I0 => sig00000c8e,
      I1 => sig00000c16,
      I2 => sig00000c32,
      O => sig00000b7a
    );
  blk000010e9 : LUT3
    generic map(
      INIT => X"D8"
    )
    port map (
      I0 => sig00000c8e,
      I1 => sig00000c18,
      I2 => sig00000c34,
      O => sig00000b78
    );
  blk000010ea : LUT3
    generic map(
      INIT => X"D8"
    )
    port map (
      I0 => sig00000c8e,
      I1 => sig00000c14,
      I2 => sig00000c30,
      O => sig00000b7c
    );
  blk000010eb : LUT3
    generic map(
      INIT => X"D8"
    )
    port map (
      I0 => sig00000c8e,
      I1 => sig00000c13,
      I2 => sig00000c2f,
      O => sig00000b7d
    );
  blk000010ec : LUT3
    generic map(
      INIT => X"D8"
    )
    port map (
      I0 => sig00000c8e,
      I1 => sig00000c15,
      I2 => sig00000c31,
      O => sig00000b7b
    );
  blk000010ed : LUT3
    generic map(
      INIT => X"D8"
    )
    port map (
      I0 => sig00000c8e,
      I1 => sig00000c12,
      I2 => sig00000c2e,
      O => sig00000b7e
    );
  blk000010ee : LUT3
    generic map(
      INIT => X"D8"
    )
    port map (
      I0 => sig00000c8e,
      I1 => sig00000c11,
      I2 => sig00000c2d,
      O => sig00000b7f
    );
  blk000010ef : LUT3
    generic map(
      INIT => X"D8"
    )
    port map (
      I0 => sig00000c8e,
      I1 => sig00000c0f,
      I2 => sig00000c2b,
      O => sig00000b81
    );
  blk000010f0 : LUT3
    generic map(
      INIT => X"D8"
    )
    port map (
      I0 => sig00000c8e,
      I1 => sig00000c38,
      I2 => sig00000c1c,
      O => sig00000b82
    );
  blk000010f1 : LUT3
    generic map(
      INIT => X"D8"
    )
    port map (
      I0 => sig00000c8e,
      I1 => sig00000c10,
      I2 => sig00000c2c,
      O => sig00000b80
    );
  blk000010f2 : LUT3
    generic map(
      INIT => X"D8"
    )
    port map (
      I0 => sig00000c8e,
      I1 => sig00000c36,
      I2 => sig00000c1a,
      O => sig00000b84
    );
  blk000010f3 : LUT3
    generic map(
      INIT => X"D8"
    )
    port map (
      I0 => sig00000c8e,
      I1 => sig00000c35,
      I2 => sig00000c19,
      O => sig00000b85
    );
  blk000010f4 : LUT3
    generic map(
      INIT => X"D8"
    )
    port map (
      I0 => sig00000c8e,
      I1 => sig00000c37,
      I2 => sig00000c1b,
      O => sig00000b83
    );
  blk000010f5 : LUT3
    generic map(
      INIT => X"D8"
    )
    port map (
      I0 => sig00000c8e,
      I1 => sig00000c33,
      I2 => sig00000c17,
      O => sig00000b87
    );
  blk000010f6 : LUT3
    generic map(
      INIT => X"D8"
    )
    port map (
      I0 => sig00000c8e,
      I1 => sig00000c32,
      I2 => sig00000c16,
      O => sig00000b88
    );
  blk000010f7 : LUT3
    generic map(
      INIT => X"D8"
    )
    port map (
      I0 => sig00000c8e,
      I1 => sig00000c34,
      I2 => sig00000c18,
      O => sig00000b86
    );
  blk000010f8 : LUT3
    generic map(
      INIT => X"D8"
    )
    port map (
      I0 => sig00000c8e,
      I1 => sig00000c31,
      I2 => sig00000c15,
      O => sig00000b89
    );
  blk000010f9 : LUT3
    generic map(
      INIT => X"D8"
    )
    port map (
      I0 => sig00000c8e,
      I1 => sig00000c30,
      I2 => sig00000c14,
      O => sig00000b8a
    );
  blk000010fa : LUT3
    generic map(
      INIT => X"D8"
    )
    port map (
      I0 => sig00000c8e,
      I1 => sig00000c2e,
      I2 => sig00000c12,
      O => sig00000b8c
    );
  blk000010fb : LUT3
    generic map(
      INIT => X"D8"
    )
    port map (
      I0 => sig00000c8e,
      I1 => sig00000c2d,
      I2 => sig00000c11,
      O => sig00000b8d
    );
  blk000010fc : LUT3
    generic map(
      INIT => X"D8"
    )
    port map (
      I0 => sig00000c8e,
      I1 => sig00000c2f,
      I2 => sig00000c13,
      O => sig00000b8b
    );
  blk000010fd : LUT3
    generic map(
      INIT => X"D8"
    )
    port map (
      I0 => sig00000c8e,
      I1 => sig00000c2b,
      I2 => sig00000c0f,
      O => sig00000b8f
    );
  blk000010fe : LUT3
    generic map(
      INIT => X"D8"
    )
    port map (
      I0 => sig00000c8e,
      I1 => sig00000c2c,
      I2 => sig00000c10,
      O => sig00000b8e
    );
  blk000010ff : LUT3
    generic map(
      INIT => X"D8"
    )
    port map (
      I0 => sig00000c90,
      I1 => sig00000c62,
      I2 => sig00000bf2,
      O => sig00000b58
    );
  blk00001100 : LUT3
    generic map(
      INIT => X"D8"
    )
    port map (
      I0 => sig00000c90,
      I1 => sig00000c61,
      I2 => sig00000bf1,
      O => sig00000b59
    );
  blk00001101 : LUT3
    generic map(
      INIT => X"D8"
    )
    port map (
      I0 => sig00000c90,
      I1 => sig00000c5f,
      I2 => sig00000bef,
      O => sig00000b5b
    );
  blk00001102 : LUT3
    generic map(
      INIT => X"D8"
    )
    port map (
      I0 => sig00000c90,
      I1 => sig00000c5e,
      I2 => sig00000bee,
      O => sig00000b5c
    );
  blk00001103 : LUT3
    generic map(
      INIT => X"D8"
    )
    port map (
      I0 => sig00000c90,
      I1 => sig00000c60,
      I2 => sig00000bf0,
      O => sig00000b5a
    );
  blk00001104 : LUT3
    generic map(
      INIT => X"D8"
    )
    port map (
      I0 => sig00000c90,
      I1 => sig00000c5d,
      I2 => sig00000bed,
      O => sig00000b5d
    );
  blk00001105 : LUT3
    generic map(
      INIT => X"D8"
    )
    port map (
      I0 => sig00000c90,
      I1 => sig00000c5c,
      I2 => sig00000bec,
      O => sig00000b5e
    );
  blk00001106 : LUT3
    generic map(
      INIT => X"D8"
    )
    port map (
      I0 => sig00000c90,
      I1 => sig00000c5a,
      I2 => sig00000bea,
      O => sig00000b60
    );
  blk00001107 : LUT3
    generic map(
      INIT => X"D8"
    )
    port map (
      I0 => sig00000c90,
      I1 => sig00000c59,
      I2 => sig00000be9,
      O => sig00000b61
    );
  blk00001108 : LUT3
    generic map(
      INIT => X"D8"
    )
    port map (
      I0 => sig00000c90,
      I1 => sig00000c5b,
      I2 => sig00000beb,
      O => sig00000b5f
    );
  blk00001109 : LUT3
    generic map(
      INIT => X"D8"
    )
    port map (
      I0 => sig00000c90,
      I1 => sig00000c57,
      I2 => sig00000be7,
      O => sig00000b63
    );
  blk0000110a : LUT3
    generic map(
      INIT => X"D8"
    )
    port map (
      I0 => sig00000c90,
      I1 => sig00000c56,
      I2 => sig00000be6,
      O => sig00000b64
    );
  blk0000110b : LUT3
    generic map(
      INIT => X"D8"
    )
    port map (
      I0 => sig00000c90,
      I1 => sig00000c58,
      I2 => sig00000be8,
      O => sig00000b62
    );
  blk0000110c : LUT3
    generic map(
      INIT => X"D8"
    )
    port map (
      I0 => sig00000c90,
      I1 => sig00000bf2,
      I2 => sig00000c62,
      O => sig00000b66
    );
  blk0000110d : LUT3
    generic map(
      INIT => X"D8"
    )
    port map (
      I0 => sig00000c90,
      I1 => sig00000bf1,
      I2 => sig00000c61,
      O => sig00000b67
    );
  blk0000110e : LUT3
    generic map(
      INIT => X"D8"
    )
    port map (
      I0 => sig00000c90,
      I1 => sig00000c55,
      I2 => sig00000be5,
      O => sig00000b65
    );
  blk0000110f : LUT3
    generic map(
      INIT => X"D8"
    )
    port map (
      I0 => sig00000c90,
      I1 => sig00000bf0,
      I2 => sig00000c60,
      O => sig00000b68
    );
  blk00001110 : LUT3
    generic map(
      INIT => X"D8"
    )
    port map (
      I0 => sig00000c90,
      I1 => sig00000bef,
      I2 => sig00000c5f,
      O => sig00000b69
    );
  blk00001111 : LUT3
    generic map(
      INIT => X"D8"
    )
    port map (
      I0 => sig00000c90,
      I1 => sig00000bed,
      I2 => sig00000c5d,
      O => sig00000b6b
    );
  blk00001112 : LUT3
    generic map(
      INIT => X"D8"
    )
    port map (
      I0 => sig00000c90,
      I1 => sig00000bec,
      I2 => sig00000c5c,
      O => sig00000b6c
    );
  blk00001113 : LUT3
    generic map(
      INIT => X"D8"
    )
    port map (
      I0 => sig00000c90,
      I1 => sig00000bee,
      I2 => sig00000c5e,
      O => sig00000b6a
    );
  blk00001114 : LUT3
    generic map(
      INIT => X"D8"
    )
    port map (
      I0 => sig00000c90,
      I1 => sig00000bea,
      I2 => sig00000c5a,
      O => sig00000b6e
    );
  blk00001115 : LUT3
    generic map(
      INIT => X"D8"
    )
    port map (
      I0 => sig00000c90,
      I1 => sig00000be9,
      I2 => sig00000c59,
      O => sig00000b6f
    );
  blk00001116 : LUT3
    generic map(
      INIT => X"D8"
    )
    port map (
      I0 => sig00000c90,
      I1 => sig00000beb,
      I2 => sig00000c5b,
      O => sig00000b6d
    );
  blk00001117 : LUT3
    generic map(
      INIT => X"D8"
    )
    port map (
      I0 => sig00000c90,
      I1 => sig00000be7,
      I2 => sig00000c57,
      O => sig00000b71
    );
  blk00001118 : LUT3
    generic map(
      INIT => X"D8"
    )
    port map (
      I0 => sig00000c90,
      I1 => sig00000be6,
      I2 => sig00000c56,
      O => sig00000b72
    );
  blk00001119 : LUT3
    generic map(
      INIT => X"D8"
    )
    port map (
      I0 => sig00000c90,
      I1 => sig00000be8,
      I2 => sig00000c58,
      O => sig00000b70
    );
  blk0000111a : LUT3
    generic map(
      INIT => X"D8"
    )
    port map (
      I0 => sig00000c90,
      I1 => sig00000be5,
      I2 => sig00000c55,
      O => sig00000b73
    );
  blk0000111b : LUT2
    generic map(
      INIT => X"8"
    )
    port map (
      I0 => sig00000c8d,
      I1 => sig00000c92,
      O => sig00000b9d
    );
  blk0000111c : LUT2
    generic map(
      INIT => X"4"
    )
    port map (
      I0 => sig00000c92,
      I1 => sig00000c8d,
      O => sig00000bc7
    );
  blk0000111d : LUT2
    generic map(
      INIT => X"8"
    )
    port map (
      I0 => sig00000a58,
      I1 => sig00000a57,
      O => sig00000be4
    );
  blk0000111e : LUT4
    generic map(
      INIT => X"EA2A"
    )
    port map (
      I0 => sig00000cc9,
      I1 => sig000000ca,
      I2 => ce,
      I3 => sig000000c9,
      O => sig00000ca9
    );
  blk0000111f : LUT3
    generic map(
      INIT => X"D8"
    )
    port map (
      I0 => ce,
      I1 => sig00000ca7,
      I2 => sig000000aa,
      O => sig00000ca8
    );
  blk00001120 : LUT3
    generic map(
      INIT => X"D8"
    )
    port map (
      I0 => sig00000d61,
      I1 => sig00000d3a,
      I2 => sig00000d54,
      O => sig00000cef
    );
  blk00001121 : LUT3
    generic map(
      INIT => X"D8"
    )
    port map (
      I0 => sig00000d61,
      I1 => sig00000d39,
      I2 => sig00000d53,
      O => sig00000cf0
    );
  blk00001122 : LUT3
    generic map(
      INIT => X"D8"
    )
    port map (
      I0 => sig00000d61,
      I1 => sig00000d38,
      I2 => sig00000d52,
      O => sig00000cf1
    );
  blk00001123 : LUT3
    generic map(
      INIT => X"D8"
    )
    port map (
      I0 => sig00000d61,
      I1 => sig00000d36,
      I2 => sig00000d50,
      O => sig00000cf3
    );
  blk00001124 : LUT3
    generic map(
      INIT => X"D8"
    )
    port map (
      I0 => sig00000d61,
      I1 => sig00000d35,
      I2 => sig00000d4f,
      O => sig00000cf4
    );
  blk00001125 : LUT3
    generic map(
      INIT => X"D8"
    )
    port map (
      I0 => sig00000d61,
      I1 => sig00000d37,
      I2 => sig00000d51,
      O => sig00000cf2
    );
  blk00001126 : LUT3
    generic map(
      INIT => X"D8"
    )
    port map (
      I0 => sig00000d61,
      I1 => sig00000d34,
      I2 => sig00000d4e,
      O => sig00000cf5
    );
  blk00001127 : LUT3
    generic map(
      INIT => X"D8"
    )
    port map (
      I0 => sig00000d61,
      I1 => sig00000d33,
      I2 => sig00000d4d,
      O => sig00000cf6
    );
  blk00001128 : LUT3
    generic map(
      INIT => X"D8"
    )
    port map (
      I0 => sig00000d61,
      I1 => sig00000d32,
      I2 => sig00000d4c,
      O => sig00000cf7
    );
  blk00001129 : LUT3
    generic map(
      INIT => X"D8"
    )
    port map (
      I0 => sig00000d61,
      I1 => sig00000d31,
      I2 => sig00000d4b,
      O => sig00000cf8
    );
  blk0000112a : LUT3
    generic map(
      INIT => X"D8"
    )
    port map (
      I0 => sig00000d61,
      I1 => sig00000d2f,
      I2 => sig00000d49,
      O => sig00000cfa
    );
  blk0000112b : LUT3
    generic map(
      INIT => X"D8"
    )
    port map (
      I0 => sig00000d61,
      I1 => sig00000d2e,
      I2 => sig00000d48,
      O => sig00000cfb
    );
  blk0000112c : LUT3
    generic map(
      INIT => X"D8"
    )
    port map (
      I0 => sig00000d61,
      I1 => sig00000d30,
      I2 => sig00000d4a,
      O => sig00000cf9
    );
  blk0000112d : LUT3
    generic map(
      INIT => X"D8"
    )
    port map (
      I0 => sig00000d61,
      I1 => sig00000d54,
      I2 => sig00000d3a,
      O => sig00000cfc
    );
  blk0000112e : LUT3
    generic map(
      INIT => X"D8"
    )
    port map (
      I0 => sig00000d61,
      I1 => sig00000d53,
      I2 => sig00000d39,
      O => sig00000cfd
    );
  blk0000112f : LUT3
    generic map(
      INIT => X"D8"
    )
    port map (
      I0 => sig00000d61,
      I1 => sig00000d52,
      I2 => sig00000d38,
      O => sig00000cfe
    );
  blk00001130 : LUT3
    generic map(
      INIT => X"D8"
    )
    port map (
      I0 => sig00000d61,
      I1 => sig00000d51,
      I2 => sig00000d37,
      O => sig00000cff
    );
  blk00001131 : LUT3
    generic map(
      INIT => X"D8"
    )
    port map (
      I0 => sig00000d61,
      I1 => sig00000d4f,
      I2 => sig00000d35,
      O => sig00000d01
    );
  blk00001132 : LUT3
    generic map(
      INIT => X"D8"
    )
    port map (
      I0 => sig00000d61,
      I1 => sig00000d4e,
      I2 => sig00000d34,
      O => sig00000d02
    );
  blk00001133 : LUT3
    generic map(
      INIT => X"D8"
    )
    port map (
      I0 => sig00000d61,
      I1 => sig00000d50,
      I2 => sig00000d36,
      O => sig00000d00
    );
  blk00001134 : LUT3
    generic map(
      INIT => X"D8"
    )
    port map (
      I0 => sig00000d61,
      I1 => sig00000d4d,
      I2 => sig00000d33,
      O => sig00000d03
    );
  blk00001135 : LUT3
    generic map(
      INIT => X"D8"
    )
    port map (
      I0 => sig00000d61,
      I1 => sig00000d4c,
      I2 => sig00000d32,
      O => sig00000d04
    );
  blk00001136 : LUT3
    generic map(
      INIT => X"D8"
    )
    port map (
      I0 => sig00000d61,
      I1 => sig00000d4b,
      I2 => sig00000d31,
      O => sig00000d05
    );
  blk00001137 : LUT3
    generic map(
      INIT => X"D8"
    )
    port map (
      I0 => sig00000d61,
      I1 => sig00000d4a,
      I2 => sig00000d30,
      O => sig00000d06
    );
  blk00001138 : LUT3
    generic map(
      INIT => X"D8"
    )
    port map (
      I0 => sig00000d61,
      I1 => sig00000d48,
      I2 => sig00000d2e,
      O => sig00000d08
    );
  blk00001139 : LUT3
    generic map(
      INIT => X"D8"
    )
    port map (
      I0 => sig00000d61,
      I1 => sig00000d49,
      I2 => sig00000d2f,
      O => sig00000d07
    );
  blk0000113a : LUT3
    generic map(
      INIT => X"D8"
    )
    port map (
      I0 => sig000000ec,
      I1 => sig00000d6f,
      I2 => sig000000e2,
      O => sig00000d09
    );
  blk0000113b : LUT3
    generic map(
      INIT => X"D8"
    )
    port map (
      I0 => sig000000ec,
      I1 => sig00000d6e,
      I2 => sig000000e1,
      O => sig00000d0a
    );
  blk0000113c : LUT3
    generic map(
      INIT => X"D8"
    )
    port map (
      I0 => sig000000ec,
      I1 => sig00000d6d,
      I2 => sig000000e0,
      O => sig00000d0b
    );
  blk0000113d : LUT3
    generic map(
      INIT => X"D8"
    )
    port map (
      I0 => sig000000ec,
      I1 => sig00000d6b,
      I2 => sig000000de,
      O => sig00000d0d
    );
  blk0000113e : LUT3
    generic map(
      INIT => X"D8"
    )
    port map (
      I0 => sig000000ec,
      I1 => sig00000d6a,
      I2 => sig000000dd,
      O => sig00000d0e
    );
  blk0000113f : LUT3
    generic map(
      INIT => X"D8"
    )
    port map (
      I0 => sig000000ec,
      I1 => sig00000d6c,
      I2 => sig000000df,
      O => sig00000d0c
    );
  blk00001140 : LUT3
    generic map(
      INIT => X"D8"
    )
    port map (
      I0 => sig000000ec,
      I1 => sig00000d69,
      I2 => sig000000dc,
      O => sig00000d0f
    );
  blk00001141 : LUT3
    generic map(
      INIT => X"D8"
    )
    port map (
      I0 => sig000000ec,
      I1 => sig00000d68,
      I2 => sig000000db,
      O => sig00000d10
    );
  blk00001142 : LUT3
    generic map(
      INIT => X"D8"
    )
    port map (
      I0 => sig000000ec,
      I1 => sig00000d67,
      I2 => sig000000da,
      O => sig00000d11
    );
  blk00001143 : LUT3
    generic map(
      INIT => X"D8"
    )
    port map (
      I0 => sig000000ec,
      I1 => sig00000d66,
      I2 => sig000000d9,
      O => sig00000d12
    );
  blk00001144 : LUT3
    generic map(
      INIT => X"D8"
    )
    port map (
      I0 => sig000000ec,
      I1 => sig00000d64,
      I2 => sig000000d7,
      O => sig00000d14
    );
  blk00001145 : LUT3
    generic map(
      INIT => X"D8"
    )
    port map (
      I0 => sig000000ec,
      I1 => sig000000e2,
      I2 => sig00000d6f,
      O => sig00000d15
    );
  blk00001146 : LUT3
    generic map(
      INIT => X"D8"
    )
    port map (
      I0 => sig000000ec,
      I1 => sig00000d65,
      I2 => sig000000d8,
      O => sig00000d13
    );
  blk00001147 : LUT3
    generic map(
      INIT => X"D8"
    )
    port map (
      I0 => sig000000ec,
      I1 => sig000000e1,
      I2 => sig00000d6e,
      O => sig00000d16
    );
  blk00001148 : LUT3
    generic map(
      INIT => X"D8"
    )
    port map (
      I0 => sig000000ec,
      I1 => sig000000e0,
      I2 => sig00000d6d,
      O => sig00000d17
    );
  blk00001149 : LUT3
    generic map(
      INIT => X"D8"
    )
    port map (
      I0 => sig000000ec,
      I1 => sig000000df,
      I2 => sig00000d6c,
      O => sig00000d18
    );
  blk0000114a : LUT3
    generic map(
      INIT => X"D8"
    )
    port map (
      I0 => sig000000ec,
      I1 => sig000000de,
      I2 => sig00000d6b,
      O => sig00000d19
    );
  blk0000114b : LUT3
    generic map(
      INIT => X"D8"
    )
    port map (
      I0 => sig000000ec,
      I1 => sig000000dd,
      I2 => sig00000d6a,
      O => sig00000d1a
    );
  blk0000114c : LUT3
    generic map(
      INIT => X"D8"
    )
    port map (
      I0 => sig000000ec,
      I1 => sig000000dc,
      I2 => sig00000d69,
      O => sig00000d1b
    );
  blk0000114d : LUT3
    generic map(
      INIT => X"D8"
    )
    port map (
      I0 => sig000000ec,
      I1 => sig000000db,
      I2 => sig00000d68,
      O => sig00000d1c
    );
  blk0000114e : LUT3
    generic map(
      INIT => X"D8"
    )
    port map (
      I0 => sig000000ec,
      I1 => sig000000da,
      I2 => sig00000d67,
      O => sig00000d1d
    );
  blk0000114f : LUT3
    generic map(
      INIT => X"D8"
    )
    port map (
      I0 => sig000000ec,
      I1 => sig000000d9,
      I2 => sig00000d66,
      O => sig00000d1e
    );
  blk00001150 : LUT3
    generic map(
      INIT => X"D8"
    )
    port map (
      I0 => sig000000ec,
      I1 => sig000000d8,
      I2 => sig00000d65,
      O => sig00000d1f
    );
  blk00001151 : LUT3
    generic map(
      INIT => X"D8"
    )
    port map (
      I0 => sig000000ec,
      I1 => sig000000d7,
      I2 => sig00000d64,
      O => sig00000d20
    );
  blk00001152 : LUT4
    generic map(
      INIT => X"7D28"
    )
    port map (
      I0 => sig00000eaf,
      I1 => sig00000ce2,
      I2 => sig00000eb4,
      I3 => sig00000cd5,
      O => sig00000dc0
    );
  blk00001153 : LUT4
    generic map(
      INIT => X"7D28"
    )
    port map (
      I0 => sig00000eaf,
      I1 => sig00000ce3,
      I2 => sig00000eb4,
      I3 => sig00000cd6,
      O => sig00000dc1
    );
  blk00001154 : LUT4
    generic map(
      INIT => X"7D28"
    )
    port map (
      I0 => sig00000eaf,
      I1 => sig00000ce5,
      I2 => sig00000eb4,
      I3 => sig00000cd8,
      O => sig00000dc3
    );
  blk00001155 : LUT4
    generic map(
      INIT => X"7D28"
    )
    port map (
      I0 => sig00000eaf,
      I1 => sig00000ce6,
      I2 => sig00000eb4,
      I3 => sig00000cd9,
      O => sig00000dc4
    );
  blk00001156 : LUT4
    generic map(
      INIT => X"7D28"
    )
    port map (
      I0 => sig00000eaf,
      I1 => sig00000ce4,
      I2 => sig00000eb4,
      I3 => sig00000cd7,
      O => sig00000dc2
    );
  blk00001157 : LUT4
    generic map(
      INIT => X"7D28"
    )
    port map (
      I0 => sig00000eaf,
      I1 => sig00000ce8,
      I2 => sig00000eb4,
      I3 => sig00000cdb,
      O => sig00000dc6
    );
  blk00001158 : LUT4
    generic map(
      INIT => X"7D28"
    )
    port map (
      I0 => sig00000eaf,
      I1 => sig00000ce9,
      I2 => sig00000eb4,
      I3 => sig00000cdc,
      O => sig00000dc7
    );
  blk00001159 : LUT4
    generic map(
      INIT => X"7D28"
    )
    port map (
      I0 => sig00000eaf,
      I1 => sig00000ce7,
      I2 => sig00000eb4,
      I3 => sig00000cda,
      O => sig00000dc5
    );
  blk0000115a : LUT4
    generic map(
      INIT => X"7D28"
    )
    port map (
      I0 => sig00000eaf,
      I1 => sig00000cea,
      I2 => sig00000eb4,
      I3 => sig00000cdd,
      O => sig00000dc8
    );
  blk0000115b : LUT4
    generic map(
      INIT => X"7D28"
    )
    port map (
      I0 => sig00000eaf,
      I1 => sig00000ceb,
      I2 => sig00000eb4,
      I3 => sig00000cde,
      O => sig00000dc9
    );
  blk0000115c : LUT4
    generic map(
      INIT => X"7D28"
    )
    port map (
      I0 => sig00000eaf,
      I1 => sig00000ced,
      I2 => sig00000eb4,
      I3 => sig00000ce0,
      O => sig00000dcb
    );
  blk0000115d : LUT4
    generic map(
      INIT => X"7D28"
    )
    port map (
      I0 => sig00000eaf,
      I1 => sig00000cee,
      I2 => sig00000eb4,
      I3 => sig00000ce1,
      O => sig00000dcc
    );
  blk0000115e : LUT4
    generic map(
      INIT => X"7D28"
    )
    port map (
      I0 => sig00000eaf,
      I1 => sig00000cec,
      I2 => sig00000eb4,
      I3 => sig00000cdf,
      O => sig00000dca
    );
  blk0000115f : LUT4
    generic map(
      INIT => X"D782"
    )
    port map (
      I0 => sig00000eaf,
      I1 => sig00000cd5,
      I2 => sig00000eb4,
      I3 => sig00000ce2,
      O => sig00000dea
    );
  blk00001160 : LUT4
    generic map(
      INIT => X"D782"
    )
    port map (
      I0 => sig00000eaf,
      I1 => sig00000cd7,
      I2 => sig00000eb4,
      I3 => sig00000ce4,
      O => sig00000dec
    );
  blk00001161 : LUT4
    generic map(
      INIT => X"D782"
    )
    port map (
      I0 => sig00000eaf,
      I1 => sig00000cd8,
      I2 => sig00000eb4,
      I3 => sig00000ce5,
      O => sig00000ded
    );
  blk00001162 : LUT4
    generic map(
      INIT => X"D782"
    )
    port map (
      I0 => sig00000eaf,
      I1 => sig00000cd6,
      I2 => sig00000eb4,
      I3 => sig00000ce3,
      O => sig00000deb
    );
  blk00001163 : LUT4
    generic map(
      INIT => X"D782"
    )
    port map (
      I0 => sig00000eaf,
      I1 => sig00000cd9,
      I2 => sig00000eb4,
      I3 => sig00000ce6,
      O => sig00000dee
    );
  blk00001164 : LUT4
    generic map(
      INIT => X"D782"
    )
    port map (
      I0 => sig00000eaf,
      I1 => sig00000cda,
      I2 => sig00000eb4,
      I3 => sig00000ce7,
      O => sig00000def
    );
  blk00001165 : LUT4
    generic map(
      INIT => X"D782"
    )
    port map (
      I0 => sig00000eaf,
      I1 => sig00000cdc,
      I2 => sig00000eb4,
      I3 => sig00000ce9,
      O => sig00000df1
    );
  blk00001166 : LUT4
    generic map(
      INIT => X"D782"
    )
    port map (
      I0 => sig00000eaf,
      I1 => sig00000cdd,
      I2 => sig00000eb4,
      I3 => sig00000cea,
      O => sig00000df2
    );
  blk00001167 : LUT4
    generic map(
      INIT => X"D782"
    )
    port map (
      I0 => sig00000eaf,
      I1 => sig00000cdb,
      I2 => sig00000eb4,
      I3 => sig00000ce8,
      O => sig00000df0
    );
  blk00001168 : LUT4
    generic map(
      INIT => X"D782"
    )
    port map (
      I0 => sig00000eaf,
      I1 => sig00000cdf,
      I2 => sig00000eb4,
      I3 => sig00000cec,
      O => sig00000df4
    );
  blk00001169 : LUT4
    generic map(
      INIT => X"D782"
    )
    port map (
      I0 => sig00000eaf,
      I1 => sig00000ce0,
      I2 => sig00000eb4,
      I3 => sig00000ced,
      O => sig00000df5
    );
  blk0000116a : LUT4
    generic map(
      INIT => X"D782"
    )
    port map (
      I0 => sig00000eaf,
      I1 => sig00000cde,
      I2 => sig00000eb4,
      I3 => sig00000ceb,
      O => sig00000df3
    );
  blk0000116b : LUT4
    generic map(
      INIT => X"D782"
    )
    port map (
      I0 => sig00000eaf,
      I1 => sig00000ce1,
      I2 => sig00000eb4,
      I3 => sig00000cee,
      O => sig00000df6
    );
  blk0000116c : LUT3
    generic map(
      INIT => X"D8"
    )
    port map (
      I0 => sig00000eb0,
      I1 => sig00000e3d,
      I2 => sig00000e59,
      O => sig00000da5
    );
  blk0000116d : LUT3
    generic map(
      INIT => X"D8"
    )
    port map (
      I0 => sig00000eb0,
      I1 => sig00000e3c,
      I2 => sig00000e58,
      O => sig00000da6
    );
  blk0000116e : LUT3
    generic map(
      INIT => X"D8"
    )
    port map (
      I0 => sig00000eb0,
      I1 => sig00000e3e,
      I2 => sig00000e5a,
      O => sig00000da4
    );
  blk0000116f : LUT3
    generic map(
      INIT => X"D8"
    )
    port map (
      I0 => sig00000eb0,
      I1 => sig00000e3b,
      I2 => sig00000e57,
      O => sig00000da7
    );
  blk00001170 : LUT3
    generic map(
      INIT => X"D8"
    )
    port map (
      I0 => sig00000eb0,
      I1 => sig00000e3a,
      I2 => sig00000e56,
      O => sig00000da8
    );
  blk00001171 : LUT3
    generic map(
      INIT => X"D8"
    )
    port map (
      I0 => sig00000eb0,
      I1 => sig00000e38,
      I2 => sig00000e54,
      O => sig00000daa
    );
  blk00001172 : LUT3
    generic map(
      INIT => X"D8"
    )
    port map (
      I0 => sig00000eb0,
      I1 => sig00000e37,
      I2 => sig00000e53,
      O => sig00000dab
    );
  blk00001173 : LUT3
    generic map(
      INIT => X"D8"
    )
    port map (
      I0 => sig00000eb0,
      I1 => sig00000e39,
      I2 => sig00000e55,
      O => sig00000da9
    );
  blk00001174 : LUT3
    generic map(
      INIT => X"D8"
    )
    port map (
      I0 => sig00000eb0,
      I1 => sig00000e35,
      I2 => sig00000e51,
      O => sig00000dad
    );
  blk00001175 : LUT3
    generic map(
      INIT => X"D8"
    )
    port map (
      I0 => sig00000eb0,
      I1 => sig00000e34,
      I2 => sig00000e50,
      O => sig00000dae
    );
  blk00001176 : LUT3
    generic map(
      INIT => X"D8"
    )
    port map (
      I0 => sig00000eb0,
      I1 => sig00000e36,
      I2 => sig00000e52,
      O => sig00000dac
    );
  blk00001177 : LUT3
    generic map(
      INIT => X"D8"
    )
    port map (
      I0 => sig00000eb0,
      I1 => sig00000e32,
      I2 => sig00000e4e,
      O => sig00000db0
    );
  blk00001178 : LUT3
    generic map(
      INIT => X"D8"
    )
    port map (
      I0 => sig00000eb0,
      I1 => sig00000e31,
      I2 => sig00000e4d,
      O => sig00000db1
    );
  blk00001179 : LUT3
    generic map(
      INIT => X"D8"
    )
    port map (
      I0 => sig00000eb0,
      I1 => sig00000e33,
      I2 => sig00000e4f,
      O => sig00000daf
    );
  blk0000117a : LUT3
    generic map(
      INIT => X"D8"
    )
    port map (
      I0 => sig00000eb0,
      I1 => sig00000e5a,
      I2 => sig00000e3e,
      O => sig00000db2
    );
  blk0000117b : LUT3
    generic map(
      INIT => X"D8"
    )
    port map (
      I0 => sig00000eb0,
      I1 => sig00000e59,
      I2 => sig00000e3d,
      O => sig00000db3
    );
  blk0000117c : LUT3
    generic map(
      INIT => X"D8"
    )
    port map (
      I0 => sig00000eb0,
      I1 => sig00000e57,
      I2 => sig00000e3b,
      O => sig00000db5
    );
  blk0000117d : LUT3
    generic map(
      INIT => X"D8"
    )
    port map (
      I0 => sig00000eb0,
      I1 => sig00000e56,
      I2 => sig00000e3a,
      O => sig00000db6
    );
  blk0000117e : LUT3
    generic map(
      INIT => X"D8"
    )
    port map (
      I0 => sig00000eb0,
      I1 => sig00000e58,
      I2 => sig00000e3c,
      O => sig00000db4
    );
  blk0000117f : LUT3
    generic map(
      INIT => X"D8"
    )
    port map (
      I0 => sig00000eb0,
      I1 => sig00000e54,
      I2 => sig00000e38,
      O => sig00000db8
    );
  blk00001180 : LUT3
    generic map(
      INIT => X"D8"
    )
    port map (
      I0 => sig00000eb0,
      I1 => sig00000e53,
      I2 => sig00000e37,
      O => sig00000db9
    );
  blk00001181 : LUT3
    generic map(
      INIT => X"D8"
    )
    port map (
      I0 => sig00000eb0,
      I1 => sig00000e55,
      I2 => sig00000e39,
      O => sig00000db7
    );
  blk00001182 : LUT3
    generic map(
      INIT => X"D8"
    )
    port map (
      I0 => sig00000eb0,
      I1 => sig00000e51,
      I2 => sig00000e35,
      O => sig00000dbb
    );
  blk00001183 : LUT3
    generic map(
      INIT => X"D8"
    )
    port map (
      I0 => sig00000eb0,
      I1 => sig00000e50,
      I2 => sig00000e34,
      O => sig00000dbc
    );
  blk00001184 : LUT3
    generic map(
      INIT => X"D8"
    )
    port map (
      I0 => sig00000eb0,
      I1 => sig00000e52,
      I2 => sig00000e36,
      O => sig00000dba
    );
  blk00001185 : LUT3
    generic map(
      INIT => X"D8"
    )
    port map (
      I0 => sig00000eb0,
      I1 => sig00000e4f,
      I2 => sig00000e33,
      O => sig00000dbd
    );
  blk00001186 : LUT3
    generic map(
      INIT => X"D8"
    )
    port map (
      I0 => sig00000eb0,
      I1 => sig00000e4e,
      I2 => sig00000e32,
      O => sig00000dbe
    );
  blk00001187 : LUT3
    generic map(
      INIT => X"D8"
    )
    port map (
      I0 => sig00000eb0,
      I1 => sig00000e4d,
      I2 => sig00000e31,
      O => sig00000dbf
    );
  blk00001188 : LUT3
    generic map(
      INIT => X"D8"
    )
    port map (
      I0 => sig00000eb2,
      I1 => sig00000e83,
      I2 => sig00000e21,
      O => sig00000d89
    );
  blk00001189 : LUT3
    generic map(
      INIT => X"D8"
    )
    port map (
      I0 => sig00000eb2,
      I1 => sig00000e82,
      I2 => sig00000e20,
      O => sig00000d8a
    );
  blk0000118a : LUT3
    generic map(
      INIT => X"D8"
    )
    port map (
      I0 => sig00000eb2,
      I1 => sig00000e84,
      I2 => sig00000e22,
      O => sig00000d88
    );
  blk0000118b : LUT3
    generic map(
      INIT => X"D8"
    )
    port map (
      I0 => sig00000eb2,
      I1 => sig00000e80,
      I2 => sig00000e1e,
      O => sig00000d8c
    );
  blk0000118c : LUT3
    generic map(
      INIT => X"D8"
    )
    port map (
      I0 => sig00000eb2,
      I1 => sig00000e7f,
      I2 => sig00000e1d,
      O => sig00000d8d
    );
  blk0000118d : LUT3
    generic map(
      INIT => X"D8"
    )
    port map (
      I0 => sig00000eb2,
      I1 => sig00000e81,
      I2 => sig00000e1f,
      O => sig00000d8b
    );
  blk0000118e : LUT3
    generic map(
      INIT => X"D8"
    )
    port map (
      I0 => sig00000eb2,
      I1 => sig00000e7d,
      I2 => sig00000e1b,
      O => sig00000d8f
    );
  blk0000118f : LUT3
    generic map(
      INIT => X"D8"
    )
    port map (
      I0 => sig00000eb2,
      I1 => sig00000e7c,
      I2 => sig00000e1a,
      O => sig00000d90
    );
  blk00001190 : LUT3
    generic map(
      INIT => X"D8"
    )
    port map (
      I0 => sig00000eb2,
      I1 => sig00000e7e,
      I2 => sig00000e1c,
      O => sig00000d8e
    );
  blk00001191 : LUT3
    generic map(
      INIT => X"D8"
    )
    port map (
      I0 => sig00000eb2,
      I1 => sig00000e7b,
      I2 => sig00000e19,
      O => sig00000d91
    );
  blk00001192 : LUT3
    generic map(
      INIT => X"D8"
    )
    port map (
      I0 => sig00000eb2,
      I1 => sig00000e7a,
      I2 => sig00000e18,
      O => sig00000d92
    );
  blk00001193 : LUT3
    generic map(
      INIT => X"D8"
    )
    port map (
      I0 => sig00000eb2,
      I1 => sig00000e78,
      I2 => sig00000e16,
      O => sig00000d94
    );
  blk00001194 : LUT3
    generic map(
      INIT => X"D8"
    )
    port map (
      I0 => sig00000eb2,
      I1 => sig00000e77,
      I2 => sig00000e15,
      O => sig00000d95
    );
  blk00001195 : LUT3
    generic map(
      INIT => X"D8"
    )
    port map (
      I0 => sig00000eb2,
      I1 => sig00000e79,
      I2 => sig00000e17,
      O => sig00000d93
    );
  blk00001196 : LUT3
    generic map(
      INIT => X"D8"
    )
    port map (
      I0 => sig00000eb2,
      I1 => sig00000e21,
      I2 => sig00000e83,
      O => sig00000d97
    );
  blk00001197 : LUT3
    generic map(
      INIT => X"D8"
    )
    port map (
      I0 => sig00000eb2,
      I1 => sig00000e20,
      I2 => sig00000e82,
      O => sig00000d98
    );
  blk00001198 : LUT3
    generic map(
      INIT => X"D8"
    )
    port map (
      I0 => sig00000eb2,
      I1 => sig00000e22,
      I2 => sig00000e84,
      O => sig00000d96
    );
  blk00001199 : LUT3
    generic map(
      INIT => X"D8"
    )
    port map (
      I0 => sig00000eb2,
      I1 => sig00000e1e,
      I2 => sig00000e80,
      O => sig00000d9a
    );
  blk0000119a : LUT3
    generic map(
      INIT => X"D8"
    )
    port map (
      I0 => sig00000eb2,
      I1 => sig00000e1d,
      I2 => sig00000e7f,
      O => sig00000d9b
    );
  blk0000119b : LUT3
    generic map(
      INIT => X"D8"
    )
    port map (
      I0 => sig00000eb2,
      I1 => sig00000e1f,
      I2 => sig00000e81,
      O => sig00000d99
    );
  blk0000119c : LUT3
    generic map(
      INIT => X"D8"
    )
    port map (
      I0 => sig00000eb2,
      I1 => sig00000e1c,
      I2 => sig00000e7e,
      O => sig00000d9c
    );
  blk0000119d : LUT3
    generic map(
      INIT => X"D8"
    )
    port map (
      I0 => sig00000eb2,
      I1 => sig00000e1b,
      I2 => sig00000e7d,
      O => sig00000d9d
    );
  blk0000119e : LUT3
    generic map(
      INIT => X"D8"
    )
    port map (
      I0 => sig00000eb2,
      I1 => sig00000e19,
      I2 => sig00000e7b,
      O => sig00000d9f
    );
  blk0000119f : LUT3
    generic map(
      INIT => X"D8"
    )
    port map (
      I0 => sig00000eb2,
      I1 => sig00000e18,
      I2 => sig00000e7a,
      O => sig00000da0
    );
  blk000011a0 : LUT3
    generic map(
      INIT => X"D8"
    )
    port map (
      I0 => sig00000eb2,
      I1 => sig00000e1a,
      I2 => sig00000e7c,
      O => sig00000d9e
    );
  blk000011a1 : LUT3
    generic map(
      INIT => X"D8"
    )
    port map (
      I0 => sig00000eb2,
      I1 => sig00000e16,
      I2 => sig00000e78,
      O => sig00000da2
    );
  blk000011a2 : LUT3
    generic map(
      INIT => X"D8"
    )
    port map (
      I0 => sig00000eb2,
      I1 => sig00000e15,
      I2 => sig00000e77,
      O => sig00000da3
    );
  blk000011a3 : LUT3
    generic map(
      INIT => X"D8"
    )
    port map (
      I0 => sig00000eb2,
      I1 => sig00000e17,
      I2 => sig00000e79,
      O => sig00000da1
    );
  blk000011a4 : LUT2
    generic map(
      INIT => X"8"
    )
    port map (
      I0 => sig00000eaf,
      I1 => sig00000eb4,
      O => sig00000dcd
    );
  blk000011a5 : LUT2
    generic map(
      INIT => X"4"
    )
    port map (
      I0 => sig00000eb4,
      I1 => sig00000eaf,
      O => sig00000df7
    );
  blk000011a6 : LUT2
    generic map(
      INIT => X"8"
    )
    port map (
      I0 => sig00000cd4,
      I1 => sig00000cd3,
      O => sig00000e14
    );
  blk000011a7 : LUT3
    generic map(
      INIT => X"D8"
    )
    port map (
      I0 => ce,
      I1 => sig00000edd,
      I2 => NlwRenamedSig_OI_xk_index(0),
      O => sig00000ed7
    );
  blk000011a8 : LUT3
    generic map(
      INIT => X"D8"
    )
    port map (
      I0 => ce,
      I1 => sig00000ede,
      I2 => NlwRenamedSig_OI_xk_index(1),
      O => sig00000ed8
    );
  blk000011a9 : LUT3
    generic map(
      INIT => X"D8"
    )
    port map (
      I0 => ce,
      I1 => sig00000edf,
      I2 => NlwRenamedSig_OI_xk_index(2),
      O => sig00000ed9
    );
  blk000011aa : LUT3
    generic map(
      INIT => X"D8"
    )
    port map (
      I0 => ce,
      I1 => sig00000ee0,
      I2 => NlwRenamedSig_OI_xk_index(3),
      O => sig00000eda
    );
  blk000011ab : LUT3
    generic map(
      INIT => X"D8"
    )
    port map (
      I0 => ce,
      I1 => sig00000ee1,
      I2 => NlwRenamedSig_OI_xk_index(4),
      O => sig00000edb
    );
  blk000011ac : LUT3
    generic map(
      INIT => X"D8"
    )
    port map (
      I0 => ce,
      I1 => sig00000ee2,
      I2 => NlwRenamedSig_OI_xk_index(5),
      O => sig00000edc
    );
  blk000011ad : LUT3
    generic map(
      INIT => X"69"
    )
    port map (
      I0 => sig00000eed,
      I1 => sig00000eea,
      I2 => sig00000eeb,
      O => sig00000ee4
    );
  blk000011ae : LUT4
    generic map(
      INIT => X"7E81"
    )
    port map (
      I0 => sig00000eed,
      I1 => sig00000eea,
      I2 => sig00000eeb,
      I3 => sig00000eec,
      O => sig00000ee3
    );
  blk000011af : LUT3
    generic map(
      INIT => X"D8"
    )
    port map (
      I0 => ce,
      I1 => sig00000ee6,
      I2 => sig00000eed,
      O => sig00000ee7
    );
  blk000011b0 : LUT3
    generic map(
      INIT => X"28"
    )
    port map (
      I0 => ce,
      I1 => NlwRenamedSig_OI_U0_i_synth_non_floating_point_arch_d_xfft_inst_done_int_d,
      I2 => sig00000eed,
      O => sig00000ee9
    );
  blk000011b1 : LUT4
    generic map(
      INIT => X"FFEF"
    )
    port map (
      I0 => sig00000eeb,
      I1 => sig00000eec,
      I2 => sig00000eea,
      I3 => sig00000eed,
      O => sig00000ee8
    );
  blk000011b2 : LUT4
    generic map(
      INIT => X"7D28"
    )
    port map (
      I0 => sig0000048e,
      I1 => sig0000027a,
      I2 => sig00000493,
      I3 => sig0000026d,
      O => sig00000eee
    );
  blk000011b3 : LUT4
    generic map(
      INIT => X"D782"
    )
    port map (
      I0 => sig0000048e,
      I1 => sig0000026d,
      I2 => sig00000493,
      I3 => sig0000027a,
      O => sig00000eef
    );
  blk000011b4 : LUT2
    generic map(
      INIT => X"6"
    )
    port map (
      I0 => sig000007f4,
      I1 => sig000007ff,
      O => sig00000ef0
    );
  blk000011b5 : LUT2
    generic map(
      INIT => X"6"
    )
    port map (
      I0 => sig00000824,
      I1 => sig000007e6,
      O => sig00000ef1
    );
  blk000011b6 : LUT2
    generic map(
      INIT => X"9"
    )
    port map (
      I0 => sig000007e6,
      I1 => sig00000824,
      O => sig00000ef2
    );
  blk000011b7 : LUT4
    generic map(
      INIT => X"7D28"
    )
    port map (
      I0 => sig00000c8d,
      I1 => sig00000a80,
      I2 => sig00000c92,
      I3 => sig00000a73,
      O => sig00000ef3
    );
  blk000011b8 : LUT4
    generic map(
      INIT => X"D782"
    )
    port map (
      I0 => sig00000c8d,
      I1 => sig00000a73,
      I2 => sig00000c92,
      I3 => sig00000a80,
      O => sig00000ef4
    );
  blk000011b9 : LUT4
    generic map(
      INIT => X"7D28"
    )
    port map (
      I0 => sig00000eaf,
      I1 => sig00000cee,
      I2 => sig00000eb4,
      I3 => sig00000ce1,
      O => sig00000ef5
    );
  blk000011ba : LUT4
    generic map(
      INIT => X"D782"
    )
    port map (
      I0 => sig00000eaf,
      I1 => sig00000ce1,
      I2 => sig00000eb4,
      I3 => sig00000cee,
      O => sig00000ef6
    );
  blk000011bb : LUT1
    generic map(
      INIT => X"2"
    )
    port map (
      I0 => sig000002ca,
      O => sig00000ef7
    );
  blk000011bc : LUT1
    generic map(
      INIT => X"2"
    )
    port map (
      I0 => sig000002cb,
      O => sig00000ef8
    );
  blk000011bd : LUT1
    generic map(
      INIT => X"2"
    )
    port map (
      I0 => sig000002cc,
      O => sig00000ef9
    );
  blk000011be : LUT1
    generic map(
      INIT => X"2"
    )
    port map (
      I0 => sig000002cd,
      O => sig00000efa
    );
  blk000011bf : LUT1
    generic map(
      INIT => X"2"
    )
    port map (
      I0 => sig000002ce,
      O => sig00000efb
    );
  blk000011c0 : LUT1
    generic map(
      INIT => X"2"
    )
    port map (
      I0 => sig000002cf,
      O => sig00000efc
    );
  blk000011c1 : LUT1
    generic map(
      INIT => X"2"
    )
    port map (
      I0 => sig000002d0,
      O => sig00000efd
    );
  blk000011c2 : LUT1
    generic map(
      INIT => X"2"
    )
    port map (
      I0 => sig000002d1,
      O => sig00000efe
    );
  blk000011c3 : LUT1
    generic map(
      INIT => X"2"
    )
    port map (
      I0 => sig000002d2,
      O => sig00000eff
    );
  blk000011c4 : LUT1
    generic map(
      INIT => X"2"
    )
    port map (
      I0 => sig000002d3,
      O => sig00000f00
    );
  blk000011c5 : LUT1
    generic map(
      INIT => X"2"
    )
    port map (
      I0 => sig000002d4,
      O => sig00000f01
    );
  blk000011c6 : LUT1
    generic map(
      INIT => X"2"
    )
    port map (
      I0 => sig000002d5,
      O => sig00000f02
    );
  blk000011c7 : LUT1
    generic map(
      INIT => X"2"
    )
    port map (
      I0 => sig000002d6,
      O => sig00000f03
    );
  blk000011c8 : LUT1
    generic map(
      INIT => X"2"
    )
    port map (
      I0 => sig000002bd,
      O => sig00000f04
    );
  blk000011c9 : LUT1
    generic map(
      INIT => X"2"
    )
    port map (
      I0 => sig000002be,
      O => sig00000f05
    );
  blk000011ca : LUT1
    generic map(
      INIT => X"2"
    )
    port map (
      I0 => sig000002bf,
      O => sig00000f06
    );
  blk000011cb : LUT1
    generic map(
      INIT => X"2"
    )
    port map (
      I0 => sig000002c0,
      O => sig00000f07
    );
  blk000011cc : LUT1
    generic map(
      INIT => X"2"
    )
    port map (
      I0 => sig000002c1,
      O => sig00000f08
    );
  blk000011cd : LUT1
    generic map(
      INIT => X"2"
    )
    port map (
      I0 => sig000002c2,
      O => sig00000f09
    );
  blk000011ce : LUT1
    generic map(
      INIT => X"2"
    )
    port map (
      I0 => sig000002c3,
      O => sig00000f0a
    );
  blk000011cf : LUT1
    generic map(
      INIT => X"2"
    )
    port map (
      I0 => sig000002c4,
      O => sig00000f0b
    );
  blk000011d0 : LUT1
    generic map(
      INIT => X"2"
    )
    port map (
      I0 => sig000002c5,
      O => sig00000f0c
    );
  blk000011d1 : LUT1
    generic map(
      INIT => X"2"
    )
    port map (
      I0 => sig000002c6,
      O => sig00000f0d
    );
  blk000011d2 : LUT1
    generic map(
      INIT => X"2"
    )
    port map (
      I0 => sig000002c7,
      O => sig00000f0e
    );
  blk000011d3 : LUT1
    generic map(
      INIT => X"2"
    )
    port map (
      I0 => sig000002c8,
      O => sig00000f0f
    );
  blk000011d4 : LUT1
    generic map(
      INIT => X"2"
    )
    port map (
      I0 => sig000002c9,
      O => sig00000f10
    );
  blk000011d5 : FDR
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      D => sig00000f11,
      R => sig000008b6,
      Q => sig00000045
    );
  blk000011d6 : FDR
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      D => sig00000f12,
      R => sig000008b6,
      Q => sig00000046
    );
  blk000011d7 : FD
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      D => sig00000f13,
      Q => sig0000018a
    );
  blk000011d8 : FD
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      D => sig00000f14,
      Q => sig00000047
    );
  blk000011d9 : LUT5
    generic map(
      INIT => X"0ACC0A0A"
    )
    port map (
      I0 => sig000000a4,
      I1 => sig000000c3,
      I2 => sig000000a2,
      I3 => sig0000005e,
      I4 => sig00000114,
      O => sig000001e0
    );
  blk000011da : LUT5
    generic map(
      INIT => X"0ACC0A0A"
    )
    port map (
      I0 => sig000000a5,
      I1 => sig000000c4,
      I2 => sig000000a2,
      I3 => sig0000005e,
      I4 => sig00000114,
      O => sig000001e1
    );
  blk000011db : LUT5
    generic map(
      INIT => X"0ACC0A0A"
    )
    port map (
      I0 => sig000000a6,
      I1 => sig000000c5,
      I2 => sig000000a2,
      I3 => sig0000005e,
      I4 => sig00000114,
      O => sig000001e2
    );
  blk000011dc : LUT5
    generic map(
      INIT => X"0ACC0A0A"
    )
    port map (
      I0 => sig000000a7,
      I1 => sig000000c6,
      I2 => sig000000a2,
      I3 => sig0000005e,
      I4 => sig00000114,
      O => sig000001e3
    );
  blk000011dd : LUT5
    generic map(
      INIT => X"0ACC0A0A"
    )
    port map (
      I0 => sig000000a8,
      I1 => sig000000c7,
      I2 => sig000000a2,
      I3 => sig0000005e,
      I4 => sig00000114,
      O => sig000001e4
    );
  blk000011de : LUT3
    generic map(
      INIT => X"75"
    )
    port map (
      I0 => sig000000a2,
      I1 => sig0000005e,
      I2 => sig00000114,
      O => sig000001df
    );
  blk000011df : LUT3
    generic map(
      INIT => X"60"
    )
    port map (
      I0 => sig00000496,
      I1 => sig00000497,
      I2 => sig0000071b,
      O => sig0000070e
    );
  blk000011e0 : LUT3
    generic map(
      INIT => X"60"
    )
    port map (
      I0 => sig00000495,
      I1 => sig00000497,
      I2 => sig00000735,
      O => sig00000728
    );
  blk000011e1 : LUT4
    generic map(
      INIT => X"BE82"
    )
    port map (
      I0 => sig0000021f,
      I1 => sig00000496,
      I2 => sig00000497,
      I3 => sig0000071a,
      O => sig0000070d
    );
  blk000011e2 : LUT4
    generic map(
      INIT => X"BE82"
    )
    port map (
      I0 => sig0000022b,
      I1 => sig00000495,
      I2 => sig00000497,
      I3 => sig00000734,
      O => sig00000727
    );
  blk000011e3 : LUT4
    generic map(
      INIT => X"BE82"
    )
    port map (
      I0 => sig0000021e,
      I1 => sig00000496,
      I2 => sig00000497,
      I3 => sig00000719,
      O => sig0000070c
    );
  blk000011e4 : LUT4
    generic map(
      INIT => X"BE82"
    )
    port map (
      I0 => sig0000022a,
      I1 => sig00000495,
      I2 => sig00000497,
      I3 => sig00000733,
      O => sig00000726
    );
  blk000011e5 : LUT3
    generic map(
      INIT => X"60"
    )
    port map (
      I0 => sig00000c94,
      I1 => sig00000c96,
      I2 => sig00000792,
      O => sig0000079d
    );
  blk000011e6 : LUT3
    generic map(
      INIT => X"60"
    )
    port map (
      I0 => sig00000c95,
      I1 => sig00000c96,
      I2 => sig000007a8,
      O => sig000007b3
    );
  blk000011e7 : LUT4
    generic map(
      INIT => X"BE82"
    )
    port map (
      I0 => sig0000021d,
      I1 => sig00000496,
      I2 => sig00000497,
      I3 => sig00000718,
      O => sig0000070b
    );
  blk000011e8 : LUT4
    generic map(
      INIT => X"BE82"
    )
    port map (
      I0 => sig00000229,
      I1 => sig00000495,
      I2 => sig00000497,
      I3 => sig00000732,
      O => sig00000725
    );
  blk000011e9 : LUT4
    generic map(
      INIT => X"BE82"
    )
    port map (
      I0 => sig00000a35,
      I1 => sig00000c94,
      I2 => sig00000c96,
      I3 => sig00000793,
      O => sig0000079e
    );
  blk000011ea : LUT4
    generic map(
      INIT => X"BE82"
    )
    port map (
      I0 => sig00000a2b,
      I1 => sig00000c95,
      I2 => sig00000c96,
      I3 => sig000007a9,
      O => sig000007b4
    );
  blk000011eb : LUT4
    generic map(
      INIT => X"BE82"
    )
    port map (
      I0 => sig0000021c,
      I1 => sig00000496,
      I2 => sig00000497,
      I3 => sig00000717,
      O => sig0000070a
    );
  blk000011ec : LUT4
    generic map(
      INIT => X"BE82"
    )
    port map (
      I0 => sig00000228,
      I1 => sig00000495,
      I2 => sig00000497,
      I3 => sig00000731,
      O => sig00000724
    );
  blk000011ed : LUT4
    generic map(
      INIT => X"BE82"
    )
    port map (
      I0 => sig00000a2f,
      I1 => sig00000c94,
      I2 => sig00000c96,
      I3 => sig00000794,
      O => sig0000079f
    );
  blk000011ee : LUT4
    generic map(
      INIT => X"BE82"
    )
    port map (
      I0 => sig00000a25,
      I1 => sig00000c95,
      I2 => sig00000c96,
      I3 => sig000007aa,
      O => sig000007b5
    );
  blk000011ef : LUT4
    generic map(
      INIT => X"BE82"
    )
    port map (
      I0 => sig0000021b,
      I1 => sig00000496,
      I2 => sig00000497,
      I3 => sig00000716,
      O => sig00000709
    );
  blk000011f0 : LUT4
    generic map(
      INIT => X"BE82"
    )
    port map (
      I0 => sig00000227,
      I1 => sig00000495,
      I2 => sig00000497,
      I3 => sig00000730,
      O => sig00000723
    );
  blk000011f1 : LUT4
    generic map(
      INIT => X"BE82"
    )
    port map (
      I0 => sig00000a29,
      I1 => sig00000c94,
      I2 => sig00000c96,
      I3 => sig00000795,
      O => sig000007a0
    );
  blk000011f2 : LUT4
    generic map(
      INIT => X"BE82"
    )
    port map (
      I0 => sig00000a29,
      I1 => sig00000c95,
      I2 => sig00000c96,
      I3 => sig000007ab,
      O => sig000007b6
    );
  blk000011f3 : LUT4
    generic map(
      INIT => X"BE82"
    )
    port map (
      I0 => sig0000021a,
      I1 => sig00000496,
      I2 => sig00000497,
      I3 => sig00000715,
      O => sig00000708
    );
  blk000011f4 : LUT4
    generic map(
      INIT => X"BE82"
    )
    port map (
      I0 => sig00000226,
      I1 => sig00000495,
      I2 => sig00000497,
      I3 => sig0000072f,
      O => sig00000722
    );
  blk000011f5 : LUT4
    generic map(
      INIT => X"BE82"
    )
    port map (
      I0 => sig00000a28,
      I1 => sig00000c94,
      I2 => sig00000c96,
      I3 => sig00000796,
      O => sig000007a1
    );
  blk000011f6 : LUT4
    generic map(
      INIT => X"BE82"
    )
    port map (
      I0 => sig00000a28,
      I1 => sig00000c95,
      I2 => sig00000c96,
      I3 => sig000007ac,
      O => sig000007b7
    );
  blk000011f7 : LUT4
    generic map(
      INIT => X"BE82"
    )
    port map (
      I0 => sig00000219,
      I1 => sig00000496,
      I2 => sig00000497,
      I3 => sig00000714,
      O => sig00000707
    );
  blk000011f8 : LUT4
    generic map(
      INIT => X"BE82"
    )
    port map (
      I0 => sig00000225,
      I1 => sig00000495,
      I2 => sig00000497,
      I3 => sig0000072e,
      O => sig00000721
    );
  blk000011f9 : LUT4
    generic map(
      INIT => X"BE82"
    )
    port map (
      I0 => sig00000a23,
      I1 => sig00000c94,
      I2 => sig00000c96,
      I3 => sig00000797,
      O => sig000007a2
    );
  blk000011fa : LUT4
    generic map(
      INIT => X"BE82"
    )
    port map (
      I0 => sig00000a23,
      I1 => sig00000c95,
      I2 => sig00000c96,
      I3 => sig000007ad,
      O => sig000007b8
    );
  blk000011fb : LUT4
    generic map(
      INIT => X"F960"
    )
    port map (
      I0 => sig00000497,
      I1 => sig00000496,
      I2 => sig00000713,
      I3 => sig00000218,
      O => sig00000706
    );
  blk000011fc : LUT4
    generic map(
      INIT => X"F960"
    )
    port map (
      I0 => sig00000497,
      I1 => sig00000495,
      I2 => sig0000072d,
      I3 => sig00000224,
      O => sig00000720
    );
  blk000011fd : LUT4
    generic map(
      INIT => X"BE82"
    )
    port map (
      I0 => sig00000a24,
      I1 => sig00000c94,
      I2 => sig00000c96,
      I3 => sig00000798,
      O => sig000007a3
    );
  blk000011fe : LUT4
    generic map(
      INIT => X"BE82"
    )
    port map (
      I0 => sig00000a22,
      I1 => sig00000c95,
      I2 => sig00000c96,
      I3 => sig000007ae,
      O => sig000007b9
    );
  blk000011ff : LUT4
    generic map(
      INIT => X"F960"
    )
    port map (
      I0 => sig00000497,
      I1 => sig00000496,
      I2 => sig00000712,
      I3 => sig00000217,
      O => sig00000705
    );
  blk00001200 : LUT4
    generic map(
      INIT => X"F960"
    )
    port map (
      I0 => sig00000497,
      I1 => sig00000495,
      I2 => sig0000072c,
      I3 => sig00000223,
      O => sig0000071f
    );
  blk00001201 : LUT4
    generic map(
      INIT => X"F960"
    )
    port map (
      I0 => sig00000c96,
      I1 => sig00000c94,
      I2 => sig00000799,
      I3 => sig00000a2f,
      O => sig000007a4
    );
  blk00001202 : LUT4
    generic map(
      INIT => X"F960"
    )
    port map (
      I0 => sig00000c96,
      I1 => sig00000c95,
      I2 => sig000007af,
      I3 => sig00000a25,
      O => sig000007ba
    );
  blk00001203 : LUT4
    generic map(
      INIT => X"F960"
    )
    port map (
      I0 => sig00000497,
      I1 => sig00000496,
      I2 => sig00000711,
      I3 => sig00000216,
      O => sig00000704
    );
  blk00001204 : LUT4
    generic map(
      INIT => X"F960"
    )
    port map (
      I0 => sig00000497,
      I1 => sig00000495,
      I2 => sig0000072b,
      I3 => sig00000222,
      O => sig0000071e
    );
  blk00001205 : LUT4
    generic map(
      INIT => X"F960"
    )
    port map (
      I0 => sig00000c96,
      I1 => sig00000c94,
      I2 => sig0000079a,
      I3 => sig00000a22,
      O => sig000007a5
    );
  blk00001206 : LUT4
    generic map(
      INIT => X"F960"
    )
    port map (
      I0 => sig00000c96,
      I1 => sig00000c95,
      I2 => sig000007b0,
      I3 => sig00000a24,
      O => sig000007bb
    );
  blk00001207 : LUT4
    generic map(
      INIT => X"F960"
    )
    port map (
      I0 => sig00000497,
      I1 => sig00000496,
      I2 => sig00000710,
      I3 => sig00000215,
      O => sig00000703
    );
  blk00001208 : LUT4
    generic map(
      INIT => X"F960"
    )
    port map (
      I0 => sig00000497,
      I1 => sig00000495,
      I2 => sig0000072a,
      I3 => sig00000221,
      O => sig0000071d
    );
  blk00001209 : LUT4
    generic map(
      INIT => X"F960"
    )
    port map (
      I0 => sig00000c96,
      I1 => sig00000c94,
      I2 => sig0000079b,
      I3 => sig00000a23,
      O => sig000007a6
    );
  blk0000120a : LUT4
    generic map(
      INIT => X"F960"
    )
    port map (
      I0 => sig00000c96,
      I1 => sig00000c95,
      I2 => sig000007b1,
      I3 => sig00000a23,
      O => sig000007bc
    );
  blk0000120b : LUT3
    generic map(
      INIT => X"6A"
    )
    port map (
      I0 => sig00000046,
      I1 => sig0000004b,
      I2 => ce,
      O => sig00000f12
    );
  blk0000120c : LUT5
    generic map(
      INIT => X"BBBF8880"
    )
    port map (
      I0 => sig00000046,
      I1 => ce,
      I2 => sig00000114,
      I3 => sig0000004a,
      I4 => sig00000045,
      O => sig00000f11
    );
  blk0000120d : LUT4
    generic map(
      INIT => X"45EF"
    )
    port map (
      I0 => sig00000060,
      I1 => sig000000a2,
      I2 => sig00000047,
      I3 => sig0000004a,
      O => sig00000f15
    );
  blk0000120e : LUT6
    generic map(
      INIT => X"7575757720202022"
    )
    port map (
      I0 => ce,
      I1 => sig0000005e,
      I2 => sig00000114,
      I3 => sig0000005f,
      I4 => sig00000f15,
      I5 => sig00000047,
      O => sig00000f14
    );
  blk0000120f : LUT4
    generic map(
      INIT => X"F960"
    )
    port map (
      I0 => sig00000497,
      I1 => sig00000496,
      I2 => sig0000070f,
      I3 => sig00000214,
      O => sig00000702
    );
  blk00001210 : LUT4
    generic map(
      INIT => X"F960"
    )
    port map (
      I0 => sig00000497,
      I1 => sig00000495,
      I2 => sig00000729,
      I3 => sig00000220,
      O => sig0000071c
    );
  blk00001211 : LUT4
    generic map(
      INIT => X"F960"
    )
    port map (
      I0 => sig00000c96,
      I1 => sig00000c94,
      I2 => sig0000079c,
      I3 => sig00000a24,
      O => sig000007a7
    );
  blk00001212 : LUT4
    generic map(
      INIT => X"F960"
    )
    port map (
      I0 => sig00000c96,
      I1 => sig00000c95,
      I2 => sig000007b2,
      I3 => sig00000a22,
      O => sig000007bd
    );
  blk00001213 : LUT4
    generic map(
      INIT => X"EA2A"
    )
    port map (
      I0 => sig0000018a,
      I1 => ce,
      I2 => fwd_inv_we,
      I3 => fwd_inv,
      O => sig00000f13
    );
  blk00001214 : LUT5
    generic map(
      INIT => X"44F44404"
    )
    port map (
      I0 => sig000000a2,
      I1 => sig000000a9,
      I2 => sig00000114,
      I3 => sig0000005e,
      I4 => sig000000c8,
      O => sig000001e5
    );
  blk00001215 : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => sig00000017,
      D => sig00000021,
      R => sig000008b6,
      Q => sig00000f16
    );
  blk00001216 : INV
    port map (
      I => sig0000021f,
      O => sig000006d3
    );
  blk00001217 : INV
    port map (
      I => sig0000021e,
      O => sig000006d5
    );
  blk00001218 : INV
    port map (
      I => sig0000021d,
      O => sig000006d7
    );
  blk00001219 : INV
    port map (
      I => sig0000021c,
      O => sig000006d9
    );
  blk0000121a : INV
    port map (
      I => sig0000021b,
      O => sig000006db
    );
  blk0000121b : INV
    port map (
      I => sig0000021a,
      O => sig000006dd
    );
  blk0000121c : INV
    port map (
      I => sig00000219,
      O => sig000006df
    );
  blk0000121d : INV
    port map (
      I => sig00000218,
      O => sig000006e1
    );
  blk0000121e : INV
    port map (
      I => sig00000217,
      O => sig000006e3
    );
  blk0000121f : INV
    port map (
      I => sig00000216,
      O => sig000006e5
    );
  blk00001220 : INV
    port map (
      I => sig00000215,
      O => sig000006e7
    );
  blk00001221 : INV
    port map (
      I => sig00000214,
      O => sig000006e9
    );
  blk00001222 : INV
    port map (
      I => sig0000022b,
      O => sig000006eb
    );
  blk00001223 : INV
    port map (
      I => sig0000022a,
      O => sig000006ed
    );
  blk00001224 : INV
    port map (
      I => sig00000229,
      O => sig000006ef
    );
  blk00001225 : INV
    port map (
      I => sig00000228,
      O => sig000006f1
    );
  blk00001226 : INV
    port map (
      I => sig00000227,
      O => sig000006f3
    );
  blk00001227 : INV
    port map (
      I => sig00000226,
      O => sig000006f5
    );
  blk00001228 : INV
    port map (
      I => sig00000225,
      O => sig000006f7
    );
  blk00001229 : INV
    port map (
      I => sig00000224,
      O => sig000006f9
    );
  blk0000122a : INV
    port map (
      I => sig00000223,
      O => sig000006fb
    );
  blk0000122b : INV
    port map (
      I => sig00000222,
      O => sig000006fd
    );
  blk0000122c : INV
    port map (
      I => sig00000221,
      O => sig000006ff
    );
  blk0000122d : INV
    port map (
      I => sig00000220,
      O => sig00000701
    );
  blk0000122e : INV
    port map (
      I => sig00000a24,
      O => sig000007be
    );
  blk0000122f : INV
    port map (
      I => sig00000a23,
      O => sig000007c0
    );
  blk00001230 : INV
    port map (
      I => sig00000a22,
      O => sig000007c2
    );
  blk00001231 : INV
    port map (
      I => sig00000a2f,
      O => sig000007c4
    );
  blk00001232 : INV
    port map (
      I => sig00000a24,
      O => sig000007c6
    );
  blk00001233 : INV
    port map (
      I => sig00000a23,
      O => sig000007c8
    );
  blk00001234 : INV
    port map (
      I => sig00000a28,
      O => sig000007ca
    );
  blk00001235 : INV
    port map (
      I => sig00000a29,
      O => sig000007cc
    );
  blk00001236 : INV
    port map (
      I => sig00000a2f,
      O => sig000007ce
    );
  blk00001237 : INV
    port map (
      I => sig00000a35,
      O => sig000007d0
    );
  blk00001238 : INV
    port map (
      I => sig00000a22,
      O => sig000007d2
    );
  blk00001239 : INV
    port map (
      I => sig00000a23,
      O => sig000007d4
    );
  blk0000123a : INV
    port map (
      I => sig00000a24,
      O => sig000007d6
    );
  blk0000123b : INV
    port map (
      I => sig00000a25,
      O => sig000007d8
    );
  blk0000123c : INV
    port map (
      I => sig00000a22,
      O => sig000007da
    );
  blk0000123d : INV
    port map (
      I => sig00000a23,
      O => sig000007dc
    );
  blk0000123e : INV
    port map (
      I => sig00000a28,
      O => sig000007de
    );
  blk0000123f : INV
    port map (
      I => sig00000a29,
      O => sig000007e0
    );
  blk00001240 : INV
    port map (
      I => sig00000a25,
      O => sig000007e2
    );
  blk00001241 : INV
    port map (
      I => sig00000a2b,
      O => sig000007e4
    );
  blk00001242 : INV
    port map (
      I => sig00000114,
      O => sig0000001a
    );
  blk00001243 : INV
    port map (
      I => sig00000198,
      O => sig00000166
    );
  blk00001244 : INV
    port map (
      I => sig00000187,
      O => sig00000171
    );
  blk00001245 : INV
    port map (
      I => sig00000188,
      O => sig00000172
    );
  blk00001246 : INV
    port map (
      I => NlwRenamedSig_OI_rfs,
      O => sig00000178
    );
  blk00001247 : INV
    port map (
      I => sig00000199,
      O => sig0000017e
    );
  blk00001248 : INV
    port map (
      I => sig0000019a,
      O => sig0000017f
    );
  blk00001249 : INV
    port map (
      I => sig0000019b,
      O => sig00000180
    );
  blk0000124a : INV
    port map (
      I => sig0000019c,
      O => sig00000181
    );
  blk0000124b : INV
    port map (
      I => sig0000019d,
      O => sig00000182
    );
  blk0000124c : INV
    port map (
      I => sig0000019e,
      O => sig00000183
    );
  blk0000124d : INV
    port map (
      I => sig000001bc,
      O => sig000001b6
    );
  blk0000124e : INV
    port map (
      I => sig000001bd,
      O => sig000001b8
    );
  blk0000124f : INV
    port map (
      I => sig000001dd,
      O => sig000001d7
    );
  blk00001250 : INV
    port map (
      I => sig000001de,
      O => sig000001d9
    );
  blk00001251 : INV
    port map (
      I => sig000002a0,
      O => sig00000298
    );
  blk00001252 : INV
    port map (
      I => sig000002b8,
      O => sig000002b0
    );
  blk00001253 : INV
    port map (
      I => sig00000aa2,
      O => sig00000a9a
    );
  blk00001254 : INV
    port map (
      I => sig00000abc,
      O => sig00000ab4
    );
  blk00001255 : INV
    port map (
      I => sig00000eea,
      O => sig00000ee5
    );
  blk00001256 : SRLC16E
    generic map(
      INIT => X"0000"
    )
    port map (
      A0 => sig000008b6,
      A1 => sig000008b6,
      A2 => sig000008b6,
      A3 => sig000008b6,
      CE => ce,
      CLK => clk,
      D => sig0000061d,
      Q => sig00000f17,
      Q15 => NLW_blk00001256_Q15_UNCONNECTED
    );
  blk00001257 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => sig00000f17,
      Q => sig00000551
    );
  blk00001258 : SRLC16E
    generic map(
      INIT => X"0000"
    )
    port map (
      A0 => sig000008b6,
      A1 => sig000008b6,
      A2 => sig000008b6,
      A3 => sig000008b6,
      CE => ce,
      CLK => clk,
      D => sig0000022c,
      Q => sig00000f18,
      Q15 => NLW_blk00001258_Q15_UNCONNECTED
    );
  blk00001259 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => sig00000f18,
      Q => sig00000494
    );
  blk0000125a : SRLC16E
    generic map(
      INIT => X"0000"
    )
    port map (
      A0 => sig000008b6,
      A1 => sig000008b6,
      A2 => sig000008b6,
      A3 => sig000008b6,
      CE => ce,
      CLK => clk,
      D => sig0000061e,
      Q => sig00000f19,
      Q15 => NLW_blk0000125a_Q15_UNCONNECTED
    );
  blk0000125b : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => sig00000f19,
      Q => sig00000550
    );
  blk0000125c : SRLC16E
    generic map(
      INIT => X"0000"
    )
    port map (
      A0 => sig000008b6,
      A1 => sig000008b6,
      A2 => sig000008b6,
      A3 => sig000008b6,
      CE => ce,
      CLK => clk,
      D => sig0000061c,
      Q => sig00000f1a,
      Q15 => NLW_blk0000125c_Q15_UNCONNECTED
    );
  blk0000125d : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => sig00000f1a,
      Q => sig00000552
    );
  blk0000125e : SRLC16E
    generic map(
      INIT => X"0000"
    )
    port map (
      A0 => sig000008b6,
      A1 => sig000008b6,
      A2 => sig000008b6,
      A3 => sig000008b6,
      CE => ce,
      CLK => clk,
      D => sig0000061b,
      Q => sig00000f1b,
      Q15 => NLW_blk0000125e_Q15_UNCONNECTED
    );
  blk0000125f : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => sig00000f1b,
      Q => sig00000553
    );
  blk00001260 : SRLC16E
    generic map(
      INIT => X"0000"
    )
    port map (
      A0 => sig000008b6,
      A1 => sig000008b6,
      A2 => sig000008b6,
      A3 => sig000008b6,
      CE => ce,
      CLK => clk,
      D => sig0000061a,
      Q => sig00000f1c,
      Q15 => NLW_blk00001260_Q15_UNCONNECTED
    );
  blk00001261 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => sig00000f1c,
      Q => sig00000554
    );
  blk00001262 : SRLC16E
    generic map(
      INIT => X"0000"
    )
    port map (
      A0 => sig000008b6,
      A1 => sig000008b6,
      A2 => sig000008b6,
      A3 => sig000008b6,
      CE => ce,
      CLK => clk,
      D => sig00000619,
      Q => sig00000f1d,
      Q15 => NLW_blk00001262_Q15_UNCONNECTED
    );
  blk00001263 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => sig00000f1d,
      Q => sig00000555
    );
  blk00001264 : SRLC16E
    generic map(
      INIT => X"0000"
    )
    port map (
      A0 => sig000008b6,
      A1 => sig000008b6,
      A2 => sig000008b6,
      A3 => sig000008b6,
      CE => ce,
      CLK => clk,
      D => sig00000618,
      Q => sig00000f1e,
      Q15 => NLW_blk00001264_Q15_UNCONNECTED
    );
  blk00001265 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => sig00000f1e,
      Q => sig00000556
    );
  blk00001266 : SRLC16E
    generic map(
      INIT => X"0000"
    )
    port map (
      A0 => sig000008b6,
      A1 => sig000008b6,
      A2 => sig000008b6,
      A3 => sig000008b6,
      CE => ce,
      CLK => clk,
      D => sig00000617,
      Q => sig00000f1f,
      Q15 => NLW_blk00001266_Q15_UNCONNECTED
    );
  blk00001267 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => sig00000f1f,
      Q => sig00000557
    );
  blk00001268 : SRLC16E
    generic map(
      INIT => X"0000"
    )
    port map (
      A0 => sig000008b6,
      A1 => sig000008b6,
      A2 => sig000008b6,
      A3 => sig000008b6,
      CE => ce,
      CLK => clk,
      D => sig00000616,
      Q => sig00000f20,
      Q15 => NLW_blk00001268_Q15_UNCONNECTED
    );
  blk00001269 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => sig00000f20,
      Q => sig00000558
    );
  blk0000126a : SRLC16E
    generic map(
      INIT => X"0000"
    )
    port map (
      A0 => sig000008b6,
      A1 => sig000008b6,
      A2 => sig000008b6,
      A3 => sig000008b6,
      CE => ce,
      CLK => clk,
      D => sig00000615,
      Q => sig00000f21,
      Q15 => NLW_blk0000126a_Q15_UNCONNECTED
    );
  blk0000126b : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => sig00000f21,
      Q => sig00000559
    );
  blk0000126c : SRLC16E
    generic map(
      INIT => X"0000"
    )
    port map (
      A0 => sig000008b6,
      A1 => sig000008b6,
      A2 => sig000008b6,
      A3 => sig000008b6,
      CE => ce,
      CLK => clk,
      D => sig00000623,
      Q => sig00000f22,
      Q15 => NLW_blk0000126c_Q15_UNCONNECTED
    );
  blk0000126d : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => sig00000f22,
      Q => sig0000055a
    );
  blk0000126e : SRLC16E
    generic map(
      INIT => X"0000"
    )
    port map (
      A0 => sig000008b6,
      A1 => sig000008b6,
      A2 => sig000008b6,
      A3 => sig000008b6,
      CE => ce,
      CLK => clk,
      D => sig0000062d,
      Q => sig00000f23,
      Q15 => NLW_blk0000126e_Q15_UNCONNECTED
    );
  blk0000126f : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => sig00000f23,
      Q => sig000005fc
    );
  blk00001270 : SRLC16E
    generic map(
      INIT => X"0000"
    )
    port map (
      A0 => sig000008b6,
      A1 => sig000008b6,
      A2 => sig000008b6,
      A3 => sig000008b6,
      CE => ce,
      CLK => clk,
      D => sig0000062c,
      Q => sig00000f24,
      Q15 => NLW_blk00001270_Q15_UNCONNECTED
    );
  blk00001271 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => sig00000f24,
      Q => sig000005fd
    );
  blk00001272 : SRLC16E
    generic map(
      INIT => X"0000"
    )
    port map (
      A0 => sig000008b6,
      A1 => sig000008b6,
      A2 => sig000008b6,
      A3 => sig000008b6,
      CE => ce,
      CLK => clk,
      D => sig0000062b,
      Q => sig00000f25,
      Q15 => NLW_blk00001272_Q15_UNCONNECTED
    );
  blk00001273 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => sig00000f25,
      Q => sig000005fe
    );
  blk00001274 : SRLC16E
    generic map(
      INIT => X"0000"
    )
    port map (
      A0 => sig000008b6,
      A1 => sig000008b6,
      A2 => sig000008b6,
      A3 => sig000008b6,
      CE => ce,
      CLK => clk,
      D => sig0000062a,
      Q => sig00000f26,
      Q15 => NLW_blk00001274_Q15_UNCONNECTED
    );
  blk00001275 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => sig00000f26,
      Q => sig000005ff
    );
  blk00001276 : SRLC16E
    generic map(
      INIT => X"0000"
    )
    port map (
      A0 => sig000008b6,
      A1 => sig000008b6,
      A2 => sig000008b6,
      A3 => sig000008b6,
      CE => ce,
      CLK => clk,
      D => sig00000629,
      Q => sig00000f27,
      Q15 => NLW_blk00001276_Q15_UNCONNECTED
    );
  blk00001277 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => sig00000f27,
      Q => sig00000600
    );
  blk00001278 : SRLC16E
    generic map(
      INIT => X"0000"
    )
    port map (
      A0 => sig000008b6,
      A1 => sig000008b6,
      A2 => sig000008b6,
      A3 => sig000008b6,
      CE => ce,
      CLK => clk,
      D => sig00000628,
      Q => sig00000f28,
      Q15 => NLW_blk00001278_Q15_UNCONNECTED
    );
  blk00001279 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => sig00000f28,
      Q => sig00000601
    );
  blk0000127a : SRLC16E
    generic map(
      INIT => X"0000"
    )
    port map (
      A0 => sig000008b6,
      A1 => sig000008b6,
      A2 => sig000008b6,
      A3 => sig000008b6,
      CE => ce,
      CLK => clk,
      D => sig00000627,
      Q => sig00000f29,
      Q15 => NLW_blk0000127a_Q15_UNCONNECTED
    );
  blk0000127b : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => sig00000f29,
      Q => sig00000602
    );
  blk0000127c : SRLC16E
    generic map(
      INIT => X"0000"
    )
    port map (
      A0 => sig000008b6,
      A1 => sig000008b6,
      A2 => sig000008b6,
      A3 => sig000008b6,
      CE => ce,
      CLK => clk,
      D => sig00000626,
      Q => sig00000f2a,
      Q15 => NLW_blk0000127c_Q15_UNCONNECTED
    );
  blk0000127d : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => sig00000f2a,
      Q => sig00000603
    );
  blk0000127e : SRLC16E
    generic map(
      INIT => X"0000"
    )
    port map (
      A0 => sig000008b6,
      A1 => sig000008b6,
      A2 => sig000008b6,
      A3 => sig000008b6,
      CE => ce,
      CLK => clk,
      D => sig00000625,
      Q => sig00000f2b,
      Q15 => NLW_blk0000127e_Q15_UNCONNECTED
    );
  blk0000127f : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => sig00000f2b,
      Q => sig00000604
    );
  blk00001280 : SRLC16E
    generic map(
      INIT => X"0000"
    )
    port map (
      A0 => sig000008b6,
      A1 => sig000008b6,
      A2 => sig000008b6,
      A3 => sig000008b6,
      CE => ce,
      CLK => clk,
      D => sig00000624,
      Q => sig00000f2c,
      Q15 => NLW_blk00001280_Q15_UNCONNECTED
    );
  blk00001281 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => sig00000f2c,
      Q => sig00000605
    );
  blk00001282 : SRLC16E
    generic map(
      INIT => X"0000"
    )
    port map (
      A0 => sig000008b6,
      A1 => sig000008b6,
      A2 => sig000008b6,
      A3 => sig000008b6,
      CE => ce,
      CLK => clk,
      D => sig000006c2,
      Q => sig00000f2d,
      Q15 => NLW_blk00001282_Q15_UNCONNECTED
    );
  blk00001283 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => sig00000f2d,
      Q => sig00000530
    );
  blk00001284 : SRLC16E
    generic map(
      INIT => X"0000"
    )
    port map (
      A0 => sig000008b6,
      A1 => sig000008b6,
      A2 => sig000008b6,
      A3 => sig000008b6,
      CE => ce,
      CLK => clk,
      D => sig000006c1,
      Q => sig00000f2e,
      Q15 => NLW_blk00001284_Q15_UNCONNECTED
    );
  blk00001285 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => sig00000f2e,
      Q => sig0000053d
    );
  blk00001286 : SRLC16E
    generic map(
      INIT => X"0000"
    )
    port map (
      A0 => sig000008b6,
      A1 => sig000008b6,
      A2 => sig000008b6,
      A3 => sig000008b6,
      CE => ce,
      CLK => clk,
      D => sig000006c0,
      Q => sig00000f2f,
      Q15 => NLW_blk00001286_Q15_UNCONNECTED
    );
  blk00001287 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => sig00000f2f,
      Q => sig0000053e
    );
  blk00001288 : SRLC16E
    generic map(
      INIT => X"0000"
    )
    port map (
      A0 => sig000008b6,
      A1 => sig000008b6,
      A2 => sig000008b6,
      A3 => sig000008b6,
      CE => ce,
      CLK => clk,
      D => sig000006bf,
      Q => sig00000f30,
      Q15 => NLW_blk00001288_Q15_UNCONNECTED
    );
  blk00001289 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => sig00000f30,
      Q => sig0000053f
    );
  blk0000128a : SRLC16E
    generic map(
      INIT => X"0000"
    )
    port map (
      A0 => sig000008b6,
      A1 => sig000008b6,
      A2 => sig000008b6,
      A3 => sig000008b6,
      CE => ce,
      CLK => clk,
      D => sig000006be,
      Q => sig00000f31,
      Q15 => NLW_blk0000128a_Q15_UNCONNECTED
    );
  blk0000128b : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => sig00000f31,
      Q => sig00000540
    );
  blk0000128c : SRLC16E
    generic map(
      INIT => X"0000"
    )
    port map (
      A0 => sig000008b6,
      A1 => sig000008b6,
      A2 => sig000008b6,
      A3 => sig000008b6,
      CE => ce,
      CLK => clk,
      D => sig000006bd,
      Q => sig00000f32,
      Q15 => NLW_blk0000128c_Q15_UNCONNECTED
    );
  blk0000128d : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => sig00000f32,
      Q => sig00000541
    );
  blk0000128e : SRLC16E
    generic map(
      INIT => X"0000"
    )
    port map (
      A0 => sig000008b6,
      A1 => sig000008b6,
      A2 => sig000008b6,
      A3 => sig000008b6,
      CE => ce,
      CLK => clk,
      D => sig000006bc,
      Q => sig00000f33,
      Q15 => NLW_blk0000128e_Q15_UNCONNECTED
    );
  blk0000128f : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => sig00000f33,
      Q => sig00000542
    );
  blk00001290 : SRLC16E
    generic map(
      INIT => X"0000"
    )
    port map (
      A0 => sig000008b6,
      A1 => sig000008b6,
      A2 => sig000008b6,
      A3 => sig000008b6,
      CE => ce,
      CLK => clk,
      D => sig000006bb,
      Q => sig00000f34,
      Q15 => NLW_blk00001290_Q15_UNCONNECTED
    );
  blk00001291 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => sig00000f34,
      Q => sig00000543
    );
  blk00001292 : SRLC16E
    generic map(
      INIT => X"0000"
    )
    port map (
      A0 => sig000008b6,
      A1 => sig000008b6,
      A2 => sig000008b6,
      A3 => sig000008b6,
      CE => ce,
      CLK => clk,
      D => sig000006ba,
      Q => sig00000f35,
      Q15 => NLW_blk00001292_Q15_UNCONNECTED
    );
  blk00001293 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => sig00000f35,
      Q => sig00000544
    );
  blk00001294 : SRLC16E
    generic map(
      INIT => X"0000"
    )
    port map (
      A0 => sig000008b6,
      A1 => sig000008b6,
      A2 => sig000008b6,
      A3 => sig000008b6,
      CE => ce,
      CLK => clk,
      D => sig000006b9,
      Q => sig00000f36,
      Q15 => NLW_blk00001294_Q15_UNCONNECTED
    );
  blk00001295 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => sig00000f36,
      Q => sig00000545
    );
  blk00001296 : SRLC16E
    generic map(
      INIT => X"0000"
    )
    port map (
      A0 => sig000008b6,
      A1 => sig000008b6,
      A2 => sig000008b6,
      A3 => sig000008b6,
      CE => ce,
      CLK => clk,
      D => sig000006b8,
      Q => sig00000f37,
      Q15 => NLW_blk00001296_Q15_UNCONNECTED
    );
  blk00001297 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => sig00000f37,
      Q => sig00000546
    );
  blk00001298 : SRLC16E
    generic map(
      INIT => X"0000"
    )
    port map (
      A0 => sig000008b6,
      A1 => sig000008b6,
      A2 => sig000008b6,
      A3 => sig000008b6,
      CE => ce,
      CLK => clk,
      D => sig000006b7,
      Q => sig00000f38,
      Q15 => NLW_blk00001298_Q15_UNCONNECTED
    );
  blk00001299 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => sig00000f38,
      Q => sig00000547
    );
  blk0000129a : SRLC16E
    generic map(
      INIT => X"0000"
    )
    port map (
      A0 => sig000008b6,
      A1 => sig000008b6,
      A2 => sig000008b6,
      A3 => sig000008b6,
      CE => ce,
      CLK => clk,
      D => sig000006b6,
      Q => sig00000f39,
      Q15 => NLW_blk0000129a_Q15_UNCONNECTED
    );
  blk0000129b : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => sig00000f39,
      Q => sig00000548
    );
  blk0000129c : SRLC16E
    generic map(
      INIT => X"0000"
    )
    port map (
      A0 => sig000008b6,
      A1 => sig000008b6,
      A2 => sig000008b6,
      A3 => sig000008b6,
      CE => ce,
      CLK => clk,
      D => sig000006b5,
      Q => sig00000f3a,
      Q15 => NLW_blk0000129c_Q15_UNCONNECTED
    );
  blk0000129d : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => sig00000f3a,
      Q => sig000005dc
    );
  blk0000129e : SRLC16E
    generic map(
      INIT => X"0000"
    )
    port map (
      A0 => sig000008b6,
      A1 => sig000008b6,
      A2 => sig000008b6,
      A3 => sig000008b6,
      CE => ce,
      CLK => clk,
      D => sig000006b4,
      Q => sig00000f3b,
      Q15 => NLW_blk0000129e_Q15_UNCONNECTED
    );
  blk0000129f : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => sig00000f3b,
      Q => sig000005e9
    );
  blk000012a0 : SRLC16E
    generic map(
      INIT => X"0000"
    )
    port map (
      A0 => sig000008b6,
      A1 => sig000008b6,
      A2 => sig000008b6,
      A3 => sig000008b6,
      CE => ce,
      CLK => clk,
      D => sig000006b3,
      Q => sig00000f3c,
      Q15 => NLW_blk000012a0_Q15_UNCONNECTED
    );
  blk000012a1 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => sig00000f3c,
      Q => sig000005ea
    );
  blk000012a2 : SRLC16E
    generic map(
      INIT => X"0000"
    )
    port map (
      A0 => sig000008b6,
      A1 => sig000008b6,
      A2 => sig000008b6,
      A3 => sig000008b6,
      CE => ce,
      CLK => clk,
      D => sig000006b2,
      Q => sig00000f3d,
      Q15 => NLW_blk000012a2_Q15_UNCONNECTED
    );
  blk000012a3 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => sig00000f3d,
      Q => sig000005eb
    );
  blk000012a4 : SRLC16E
    generic map(
      INIT => X"0000"
    )
    port map (
      A0 => sig000008b6,
      A1 => sig000008b6,
      A2 => sig000008b6,
      A3 => sig000008b6,
      CE => ce,
      CLK => clk,
      D => sig000006b1,
      Q => sig00000f3e,
      Q15 => NLW_blk000012a4_Q15_UNCONNECTED
    );
  blk000012a5 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => sig00000f3e,
      Q => sig000005ec
    );
  blk000012a6 : SRLC16E
    generic map(
      INIT => X"0000"
    )
    port map (
      A0 => sig000008b6,
      A1 => sig000008b6,
      A2 => sig000008b6,
      A3 => sig000008b6,
      CE => ce,
      CLK => clk,
      D => sig000006b0,
      Q => sig00000f3f,
      Q15 => NLW_blk000012a6_Q15_UNCONNECTED
    );
  blk000012a7 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => sig00000f3f,
      Q => sig000005ed
    );
  blk000012a8 : SRLC16E
    generic map(
      INIT => X"0000"
    )
    port map (
      A0 => sig000008b6,
      A1 => sig000008b6,
      A2 => sig000008b6,
      A3 => sig000008b6,
      CE => ce,
      CLK => clk,
      D => sig000006af,
      Q => sig00000f40,
      Q15 => NLW_blk000012a8_Q15_UNCONNECTED
    );
  blk000012a9 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => sig00000f40,
      Q => sig000005ee
    );
  blk000012aa : SRLC16E
    generic map(
      INIT => X"0000"
    )
    port map (
      A0 => sig000008b6,
      A1 => sig000008b6,
      A2 => sig000008b6,
      A3 => sig000008b6,
      CE => ce,
      CLK => clk,
      D => sig000006ae,
      Q => sig00000f41,
      Q15 => NLW_blk000012aa_Q15_UNCONNECTED
    );
  blk000012ab : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => sig00000f41,
      Q => sig000005ef
    );
  blk000012ac : SRLC16E
    generic map(
      INIT => X"0000"
    )
    port map (
      A0 => sig000008b6,
      A1 => sig000008b6,
      A2 => sig000008b6,
      A3 => sig000008b6,
      CE => ce,
      CLK => clk,
      D => sig000006ad,
      Q => sig00000f42,
      Q15 => NLW_blk000012ac_Q15_UNCONNECTED
    );
  blk000012ad : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => sig00000f42,
      Q => sig000005f0
    );
  blk000012ae : SRLC16E
    generic map(
      INIT => X"0000"
    )
    port map (
      A0 => sig000008b6,
      A1 => sig000008b6,
      A2 => sig000008b6,
      A3 => sig000008b6,
      CE => ce,
      CLK => clk,
      D => sig000006ac,
      Q => sig00000f43,
      Q15 => NLW_blk000012ae_Q15_UNCONNECTED
    );
  blk000012af : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => sig00000f43,
      Q => sig000005f1
    );
  blk000012b0 : SRLC16E
    generic map(
      INIT => X"0000"
    )
    port map (
      A0 => sig000008b6,
      A1 => sig000008b6,
      A2 => sig000008b6,
      A3 => sig000008b6,
      CE => ce,
      CLK => clk,
      D => sig000006ab,
      Q => sig00000f44,
      Q15 => NLW_blk000012b0_Q15_UNCONNECTED
    );
  blk000012b1 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => sig00000f44,
      Q => sig000005f2
    );
  blk000012b2 : SRLC16E
    generic map(
      INIT => X"0000"
    )
    port map (
      A0 => sig000008b6,
      A1 => sig000008b6,
      A2 => sig000008b6,
      A3 => sig000008b6,
      CE => ce,
      CLK => clk,
      D => sig000006aa,
      Q => sig00000f45,
      Q15 => NLW_blk000012b2_Q15_UNCONNECTED
    );
  blk000012b3 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => sig00000f45,
      Q => sig000005f3
    );
  blk000012b4 : SRLC16E
    generic map(
      INIT => X"0000"
    )
    port map (
      A0 => sig000008b6,
      A1 => sig000008b6,
      A2 => sig000008b6,
      A3 => sig000008b6,
      CE => ce,
      CLK => clk,
      D => sig000006a9,
      Q => sig00000f46,
      Q15 => NLW_blk000012b4_Q15_UNCONNECTED
    );
  blk000012b5 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => sig00000f46,
      Q => sig000005f4
    );
  blk000012b6 : SRLC16E
    generic map(
      INIT => X"0000"
    )
    port map (
      A0 => sig000008b6,
      A1 => sig000008b6,
      A2 => sig000008b6,
      A3 => sig000008b6,
      CE => ce,
      CLK => clk,
      D => sig00000809,
      Q => sig00000f47,
      Q15 => NLW_blk000012b6_Q15_UNCONNECTED
    );
  blk000012b7 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => sig00000f47,
      Q => sig00000823
    );
  blk000012b8 : SRLC16E
    generic map(
      INIT => X"0000"
    )
    port map (
      A0 => sig000008b6,
      A1 => sig000008b6,
      A2 => sig000008b6,
      A3 => sig000008b6,
      CE => ce,
      CLK => clk,
      D => sig00000808,
      Q => sig00000f48,
      Q15 => NLW_blk000012b8_Q15_UNCONNECTED
    );
  blk000012b9 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => sig00000f48,
      Q => sig00000822
    );
  blk000012ba : SRLC16E
    generic map(
      INIT => X"0000"
    )
    port map (
      A0 => sig000008b6,
      A1 => sig000008b6,
      A2 => sig000008b6,
      A3 => sig000008b6,
      CE => ce,
      CLK => clk,
      D => sig00000807,
      Q => sig00000f49,
      Q15 => NLW_blk000012ba_Q15_UNCONNECTED
    );
  blk000012bb : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => sig00000f49,
      Q => sig00000821
    );
  blk000012bc : SRLC16E
    generic map(
      INIT => X"0000"
    )
    port map (
      A0 => sig000008b6,
      A1 => sig000008b6,
      A2 => sig000008b6,
      A3 => sig000008b6,
      CE => ce,
      CLK => clk,
      D => sig00000806,
      Q => sig00000f4a,
      Q15 => NLW_blk000012bc_Q15_UNCONNECTED
    );
  blk000012bd : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => sig00000f4a,
      Q => sig00000820
    );
  blk000012be : SRLC16E
    generic map(
      INIT => X"0000"
    )
    port map (
      A0 => sig000008b6,
      A1 => sig000008b6,
      A2 => sig000008b6,
      A3 => sig000008b6,
      CE => ce,
      CLK => clk,
      D => sig00000805,
      Q => sig00000f4b,
      Q15 => NLW_blk000012be_Q15_UNCONNECTED
    );
  blk000012bf : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => sig00000f4b,
      Q => sig0000081f
    );
  blk000012c0 : SRLC16E
    generic map(
      INIT => X"0000"
    )
    port map (
      A0 => sig000008b6,
      A1 => sig000008b6,
      A2 => sig000008b6,
      A3 => sig000008b6,
      CE => ce,
      CLK => clk,
      D => sig00000804,
      Q => sig00000f4c,
      Q15 => NLW_blk000012c0_Q15_UNCONNECTED
    );
  blk000012c1 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => sig00000f4c,
      Q => sig0000081e
    );
  blk000012c2 : SRLC16E
    generic map(
      INIT => X"0000"
    )
    port map (
      A0 => sig000008b6,
      A1 => sig000008b6,
      A2 => sig000008b6,
      A3 => sig000008b6,
      CE => ce,
      CLK => clk,
      D => sig00000803,
      Q => sig00000f4d,
      Q15 => NLW_blk000012c2_Q15_UNCONNECTED
    );
  blk000012c3 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => sig00000f4d,
      Q => sig0000081d
    );
  blk000012c4 : SRLC16E
    generic map(
      INIT => X"0000"
    )
    port map (
      A0 => sig000008b6,
      A1 => sig000008b6,
      A2 => sig000008b6,
      A3 => sig000008b6,
      CE => ce,
      CLK => clk,
      D => sig00000802,
      Q => sig00000f4e,
      Q15 => NLW_blk000012c4_Q15_UNCONNECTED
    );
  blk000012c5 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => sig00000f4e,
      Q => sig0000081c
    );
  blk000012c6 : SRLC16E
    generic map(
      INIT => X"0000"
    )
    port map (
      A0 => sig000008b6,
      A1 => sig000008b6,
      A2 => sig000008b6,
      A3 => sig000008b6,
      CE => ce,
      CLK => clk,
      D => sig00000801,
      Q => sig00000f4f,
      Q15 => NLW_blk000012c6_Q15_UNCONNECTED
    );
  blk000012c7 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => sig00000f4f,
      Q => sig0000081b
    );
  blk000012c8 : SRLC16E
    generic map(
      INIT => X"0000"
    )
    port map (
      A0 => sig000008b6,
      A1 => sig000008b6,
      A2 => sig000008b6,
      A3 => sig000008b6,
      CE => ce,
      CLK => clk,
      D => sig00000800,
      Q => sig00000f50,
      Q15 => NLW_blk000012c8_Q15_UNCONNECTED
    );
  blk000012c9 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => sig00000f50,
      Q => sig0000081a
    );
  blk000012ca : SRLC16E
    generic map(
      INIT => X"0000"
    )
    port map (
      A0 => sig000008b6,
      A1 => sig000008b6,
      A2 => sig000008b6,
      A3 => sig000008b6,
      CE => ce,
      CLK => clk,
      D => sig000007ff,
      Q => sig00000f51,
      Q15 => NLW_blk000012ca_Q15_UNCONNECTED
    );
  blk000012cb : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => sig00000f51,
      Q => sig00000819
    );
  blk000012cc : SRLC16E
    generic map(
      INIT => X"0000"
    )
    port map (
      A0 => sig000008b6,
      A1 => sig000008b6,
      A2 => sig000008b6,
      A3 => sig000008b6,
      CE => ce,
      CLK => clk,
      D => sig000007fe,
      Q => sig00000f52,
      Q15 => NLW_blk000012cc_Q15_UNCONNECTED
    );
  blk000012cd : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => sig00000f52,
      Q => sig00000866
    );
  blk000012ce : SRLC16E
    generic map(
      INIT => X"0000"
    )
    port map (
      A0 => sig000008b6,
      A1 => sig000008b6,
      A2 => sig000008b6,
      A3 => sig000008b6,
      CE => ce,
      CLK => clk,
      D => sig000007fd,
      Q => sig00000f53,
      Q15 => NLW_blk000012ce_Q15_UNCONNECTED
    );
  blk000012cf : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => sig00000f53,
      Q => sig00000865
    );
  blk000012d0 : SRLC16E
    generic map(
      INIT => X"0000"
    )
    port map (
      A0 => sig000008b6,
      A1 => sig000008b6,
      A2 => sig000008b6,
      A3 => sig000008b6,
      CE => ce,
      CLK => clk,
      D => sig000007fc,
      Q => sig00000f54,
      Q15 => NLW_blk000012d0_Q15_UNCONNECTED
    );
  blk000012d1 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => sig00000f54,
      Q => sig00000864
    );
  blk000012d2 : SRLC16E
    generic map(
      INIT => X"0000"
    )
    port map (
      A0 => sig000008b6,
      A1 => sig000008b6,
      A2 => sig000008b6,
      A3 => sig000008b6,
      CE => ce,
      CLK => clk,
      D => sig000007fb,
      Q => sig00000f55,
      Q15 => NLW_blk000012d2_Q15_UNCONNECTED
    );
  blk000012d3 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => sig00000f55,
      Q => sig00000863
    );
  blk000012d4 : SRLC16E
    generic map(
      INIT => X"0000"
    )
    port map (
      A0 => sig000008b6,
      A1 => sig000008b6,
      A2 => sig000008b6,
      A3 => sig000008b6,
      CE => ce,
      CLK => clk,
      D => sig000007fa,
      Q => sig00000f56,
      Q15 => NLW_blk000012d4_Q15_UNCONNECTED
    );
  blk000012d5 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => sig00000f56,
      Q => sig00000862
    );
  blk000012d6 : SRLC16E
    generic map(
      INIT => X"0000"
    )
    port map (
      A0 => sig000008b6,
      A1 => sig000008b6,
      A2 => sig000008b6,
      A3 => sig000008b6,
      CE => ce,
      CLK => clk,
      D => sig000007f9,
      Q => sig00000f57,
      Q15 => NLW_blk000012d6_Q15_UNCONNECTED
    );
  blk000012d7 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => sig00000f57,
      Q => sig00000861
    );
  blk000012d8 : SRLC16E
    generic map(
      INIT => X"0000"
    )
    port map (
      A0 => sig000008b6,
      A1 => sig000008b6,
      A2 => sig000008b6,
      A3 => sig000008b6,
      CE => ce,
      CLK => clk,
      D => sig000007f6,
      Q => sig00000f58,
      Q15 => NLW_blk000012d8_Q15_UNCONNECTED
    );
  blk000012d9 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => sig00000f58,
      Q => sig0000085e
    );
  blk000012da : SRLC16E
    generic map(
      INIT => X"0000"
    )
    port map (
      A0 => sig000008b6,
      A1 => sig000008b6,
      A2 => sig000008b6,
      A3 => sig000008b6,
      CE => ce,
      CLK => clk,
      D => sig000007f8,
      Q => sig00000f59,
      Q15 => NLW_blk000012da_Q15_UNCONNECTED
    );
  blk000012db : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => sig00000f59,
      Q => sig00000860
    );
  blk000012dc : SRLC16E
    generic map(
      INIT => X"0000"
    )
    port map (
      A0 => sig000008b6,
      A1 => sig000008b6,
      A2 => sig000008b6,
      A3 => sig000008b6,
      CE => ce,
      CLK => clk,
      D => sig000007f7,
      Q => sig00000f5a,
      Q15 => NLW_blk000012dc_Q15_UNCONNECTED
    );
  blk000012dd : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => sig00000f5a,
      Q => sig0000085f
    );
  blk000012de : SRLC16E
    generic map(
      INIT => X"0000"
    )
    port map (
      A0 => sig000008b6,
      A1 => sig000008b6,
      A2 => sig000008b6,
      A3 => sig000008b6,
      CE => ce,
      CLK => clk,
      D => sig000007f5,
      Q => sig00000f5b,
      Q15 => NLW_blk000012de_Q15_UNCONNECTED
    );
  blk000012df : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => sig00000f5b,
      Q => sig0000085d
    );
  blk000012e0 : SRLC16E
    generic map(
      INIT => X"0000"
    )
    port map (
      A0 => sig000008b6,
      A1 => sig000008b6,
      A2 => sig000008b6,
      A3 => sig000008b6,
      CE => ce,
      CLK => clk,
      D => sig000007f4,
      Q => sig00000f5c,
      Q15 => NLW_blk000012e0_Q15_UNCONNECTED
    );
  blk000012e1 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => sig00000f5c,
      Q => sig0000085c
    );
  blk000012e2 : SRLC16E
    generic map(
      INIT => X"0000"
    )
    port map (
      A0 => sig000008b6,
      A1 => sig000008b6,
      A2 => sig000008b6,
      A3 => sig000008b6,
      CE => ce,
      CLK => clk,
      D => sig00000897,
      Q => sig00000f5d,
      Q15 => NLW_blk000012e2_Q15_UNCONNECTED
    );
  blk000012e3 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => sig00000f5d,
      Q => sig00000818
    );
  blk000012e4 : SRLC16E
    generic map(
      INIT => X"0000"
    )
    port map (
      A0 => sig000008b6,
      A1 => sig000008b6,
      A2 => sig000008b6,
      A3 => sig000008b6,
      CE => ce,
      CLK => clk,
      D => sig00000888,
      Q => sig00000f5e,
      Q15 => NLW_blk000012e4_Q15_UNCONNECTED
    );
  blk000012e5 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => sig00000f5e,
      Q => sig00000817
    );
  blk000012e6 : SRLC16E
    generic map(
      INIT => X"0000"
    )
    port map (
      A0 => sig000008b6,
      A1 => sig000008b6,
      A2 => sig000008b6,
      A3 => sig000008b6,
      CE => ce,
      CLK => clk,
      D => sig00000887,
      Q => sig00000f5f,
      Q15 => NLW_blk000012e6_Q15_UNCONNECTED
    );
  blk000012e7 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => sig00000f5f,
      Q => sig00000816
    );
  blk000012e8 : SRLC16E
    generic map(
      INIT => X"0000"
    )
    port map (
      A0 => sig000008b6,
      A1 => sig000008b6,
      A2 => sig000008b6,
      A3 => sig000008b6,
      CE => ce,
      CLK => clk,
      D => sig00000886,
      Q => sig00000f60,
      Q15 => NLW_blk000012e8_Q15_UNCONNECTED
    );
  blk000012e9 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => sig00000f60,
      Q => sig00000815
    );
  blk000012ea : SRLC16E
    generic map(
      INIT => X"0000"
    )
    port map (
      A0 => sig000008b6,
      A1 => sig000008b6,
      A2 => sig000008b6,
      A3 => sig000008b6,
      CE => ce,
      CLK => clk,
      D => sig00000885,
      Q => sig00000f61,
      Q15 => NLW_blk000012ea_Q15_UNCONNECTED
    );
  blk000012eb : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => sig00000f61,
      Q => sig00000814
    );
  blk000012ec : SRLC16E
    generic map(
      INIT => X"0000"
    )
    port map (
      A0 => sig000008b6,
      A1 => sig000008b6,
      A2 => sig000008b6,
      A3 => sig000008b6,
      CE => ce,
      CLK => clk,
      D => sig00000884,
      Q => sig00000f62,
      Q15 => NLW_blk000012ec_Q15_UNCONNECTED
    );
  blk000012ed : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => sig00000f62,
      Q => sig00000813
    );
  blk000012ee : SRLC16E
    generic map(
      INIT => X"0000"
    )
    port map (
      A0 => sig000008b6,
      A1 => sig000008b6,
      A2 => sig000008b6,
      A3 => sig000008b6,
      CE => ce,
      CLK => clk,
      D => sig00000883,
      Q => sig00000f63,
      Q15 => NLW_blk000012ee_Q15_UNCONNECTED
    );
  blk000012ef : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => sig00000f63,
      Q => sig00000812
    );
  blk000012f0 : SRLC16E
    generic map(
      INIT => X"0000"
    )
    port map (
      A0 => sig000008b6,
      A1 => sig000008b6,
      A2 => sig000008b6,
      A3 => sig000008b6,
      CE => ce,
      CLK => clk,
      D => sig00000882,
      Q => sig00000f64,
      Q15 => NLW_blk000012f0_Q15_UNCONNECTED
    );
  blk000012f1 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => sig00000f64,
      Q => sig00000811
    );
  blk000012f2 : SRLC16E
    generic map(
      INIT => X"0000"
    )
    port map (
      A0 => sig000008b6,
      A1 => sig000008b6,
      A2 => sig000008b6,
      A3 => sig000008b6,
      CE => ce,
      CLK => clk,
      D => sig00000881,
      Q => sig00000f65,
      Q15 => NLW_blk000012f2_Q15_UNCONNECTED
    );
  blk000012f3 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => sig00000f65,
      Q => sig00000810
    );
  blk000012f4 : SRLC16E
    generic map(
      INIT => X"0000"
    )
    port map (
      A0 => sig000008b6,
      A1 => sig000008b6,
      A2 => sig000008b6,
      A3 => sig000008b6,
      CE => ce,
      CLK => clk,
      D => sig00000880,
      Q => sig00000f66,
      Q15 => NLW_blk000012f4_Q15_UNCONNECTED
    );
  blk000012f5 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => sig00000f66,
      Q => sig0000080f
    );
  blk000012f6 : SRLC16E
    generic map(
      INIT => X"0000"
    )
    port map (
      A0 => sig000008b6,
      A1 => sig000008b6,
      A2 => sig000008b6,
      A3 => sig000008b6,
      CE => ce,
      CLK => clk,
      D => sig0000087f,
      Q => sig00000f67,
      Q15 => NLW_blk000012f6_Q15_UNCONNECTED
    );
  blk000012f7 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => sig00000f67,
      Q => sig0000080e
    );
  blk000012f8 : SRLC16E
    generic map(
      INIT => X"0000"
    )
    port map (
      A0 => sig000008b6,
      A1 => sig000008b6,
      A2 => sig000008b6,
      A3 => sig000008b6,
      CE => ce,
      CLK => clk,
      D => sig00000896,
      Q => sig00000f68,
      Q15 => NLW_blk000012f8_Q15_UNCONNECTED
    );
  blk000012f9 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => sig00000f68,
      Q => sig0000085b
    );
  blk000012fa : SRLC16E
    generic map(
      INIT => X"0000"
    )
    port map (
      A0 => sig000008b6,
      A1 => sig000008b6,
      A2 => sig000008b6,
      A3 => sig000008b6,
      CE => ce,
      CLK => clk,
      D => sig00000895,
      Q => sig00000f69,
      Q15 => NLW_blk000012fa_Q15_UNCONNECTED
    );
  blk000012fb : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => sig00000f69,
      Q => sig0000085a
    );
  blk000012fc : SRLC16E
    generic map(
      INIT => X"0000"
    )
    port map (
      A0 => sig000008b6,
      A1 => sig000008b6,
      A2 => sig000008b6,
      A3 => sig000008b6,
      CE => ce,
      CLK => clk,
      D => sig00000894,
      Q => sig00000f6a,
      Q15 => NLW_blk000012fc_Q15_UNCONNECTED
    );
  blk000012fd : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => sig00000f6a,
      Q => sig00000859
    );
  blk000012fe : SRLC16E
    generic map(
      INIT => X"0000"
    )
    port map (
      A0 => sig000008b6,
      A1 => sig000008b6,
      A2 => sig000008b6,
      A3 => sig000008b6,
      CE => ce,
      CLK => clk,
      D => sig00000893,
      Q => sig00000f6b,
      Q15 => NLW_blk000012fe_Q15_UNCONNECTED
    );
  blk000012ff : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => sig00000f6b,
      Q => sig00000858
    );
  blk00001300 : SRLC16E
    generic map(
      INIT => X"0000"
    )
    port map (
      A0 => sig000008b6,
      A1 => sig000008b6,
      A2 => sig000008b6,
      A3 => sig000008b6,
      CE => ce,
      CLK => clk,
      D => sig00000892,
      Q => sig00000f6c,
      Q15 => NLW_blk00001300_Q15_UNCONNECTED
    );
  blk00001301 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => sig00000f6c,
      Q => sig00000857
    );
  blk00001302 : SRLC16E
    generic map(
      INIT => X"0000"
    )
    port map (
      A0 => sig000008b6,
      A1 => sig000008b6,
      A2 => sig000008b6,
      A3 => sig000008b6,
      CE => ce,
      CLK => clk,
      D => sig00000891,
      Q => sig00000f6d,
      Q15 => NLW_blk00001302_Q15_UNCONNECTED
    );
  blk00001303 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => sig00000f6d,
      Q => sig00000856
    );
  blk00001304 : SRLC16E
    generic map(
      INIT => X"0000"
    )
    port map (
      A0 => sig000008b6,
      A1 => sig000008b6,
      A2 => sig000008b6,
      A3 => sig000008b6,
      CE => ce,
      CLK => clk,
      D => sig00000890,
      Q => sig00000f6e,
      Q15 => NLW_blk00001304_Q15_UNCONNECTED
    );
  blk00001305 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => sig00000f6e,
      Q => sig00000855
    );
  blk00001306 : SRLC16E
    generic map(
      INIT => X"0000"
    )
    port map (
      A0 => sig000008b6,
      A1 => sig000008b6,
      A2 => sig000008b6,
      A3 => sig000008b6,
      CE => ce,
      CLK => clk,
      D => sig0000088f,
      Q => sig00000f6f,
      Q15 => NLW_blk00001306_Q15_UNCONNECTED
    );
  blk00001307 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => sig00000f6f,
      Q => sig00000854
    );
  blk00001308 : SRLC16E
    generic map(
      INIT => X"0000"
    )
    port map (
      A0 => sig000008b6,
      A1 => sig000008b6,
      A2 => sig000008b6,
      A3 => sig000008b6,
      CE => ce,
      CLK => clk,
      D => sig0000088e,
      Q => sig00000f70,
      Q15 => NLW_blk00001308_Q15_UNCONNECTED
    );
  blk00001309 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => sig00000f70,
      Q => sig00000853
    );
  blk0000130a : SRLC16E
    generic map(
      INIT => X"0000"
    )
    port map (
      A0 => sig000008b6,
      A1 => sig000008b6,
      A2 => sig000008b6,
      A3 => sig000008b6,
      CE => ce,
      CLK => clk,
      D => sig0000088d,
      Q => sig00000f71,
      Q15 => NLW_blk0000130a_Q15_UNCONNECTED
    );
  blk0000130b : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => sig00000f71,
      Q => sig00000852
    );
  blk0000130c : SRLC16E
    generic map(
      INIT => X"0000"
    )
    port map (
      A0 => sig000008b6,
      A1 => sig000008b6,
      A2 => sig000008b6,
      A3 => sig000008b6,
      CE => ce,
      CLK => clk,
      D => sig00000a36,
      Q => sig00000f72,
      Q15 => NLW_blk0000130c_Q15_UNCONNECTED
    );
  blk0000130d : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => sig00000f72,
      Q => sig00000c93
    );
  blk0000130e : SRLC16E
    generic map(
      INIT => X"0000"
    )
    port map (
      A0 => sig000008b6,
      A1 => sig000008b6,
      A2 => sig000008b6,
      A3 => sig000008b6,
      CE => ce,
      CLK => clk,
      D => sig00000ea0,
      Q => sig00000f73,
      Q15 => NLW_blk0000130e_Q15_UNCONNECTED
    );
  blk0000130f : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => sig00000f73,
      Q => sig00000e84
    );
  blk00001310 : SRLC16E
    generic map(
      INIT => X"0000"
    )
    port map (
      A0 => sig000008b6,
      A1 => sig000008b6,
      A2 => sig000008b6,
      A3 => sig000008b6,
      CE => ce,
      CLK => clk,
      D => sig00000e9f,
      Q => sig00000f74,
      Q15 => NLW_blk00001310_Q15_UNCONNECTED
    );
  blk00001311 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => sig00000f74,
      Q => sig00000e83
    );
  blk00001312 : SRLC16E
    generic map(
      INIT => X"0000"
    )
    port map (
      A0 => sig000008b6,
      A1 => sig000008b6,
      A2 => sig000008b6,
      A3 => sig000008b6,
      CE => ce,
      CLK => clk,
      D => sig00000e9e,
      Q => sig00000f75,
      Q15 => NLW_blk00001312_Q15_UNCONNECTED
    );
  blk00001313 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => sig00000f75,
      Q => sig00000e82
    );
  blk00001314 : SRLC16E
    generic map(
      INIT => X"0000"
    )
    port map (
      A0 => sig000008b6,
      A1 => sig000008b6,
      A2 => sig000008b6,
      A3 => sig000008b6,
      CE => ce,
      CLK => clk,
      D => sig00000e9d,
      Q => sig00000f76,
      Q15 => NLW_blk00001314_Q15_UNCONNECTED
    );
  blk00001315 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => sig00000f76,
      Q => sig00000e81
    );
  blk00001316 : SRLC16E
    generic map(
      INIT => X"0000"
    )
    port map (
      A0 => sig000008b6,
      A1 => sig000008b6,
      A2 => sig000008b6,
      A3 => sig000008b6,
      CE => ce,
      CLK => clk,
      D => sig00000e9c,
      Q => sig00000f77,
      Q15 => NLW_blk00001316_Q15_UNCONNECTED
    );
  blk00001317 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => sig00000f77,
      Q => sig00000e80
    );
  blk00001318 : SRLC16E
    generic map(
      INIT => X"0000"
    )
    port map (
      A0 => sig000008b6,
      A1 => sig000008b6,
      A2 => sig000008b6,
      A3 => sig000008b6,
      CE => ce,
      CLK => clk,
      D => sig00000e9b,
      Q => sig00000f78,
      Q15 => NLW_blk00001318_Q15_UNCONNECTED
    );
  blk00001319 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => sig00000f78,
      Q => sig00000e7f
    );
  blk0000131a : SRLC16E
    generic map(
      INIT => X"0000"
    )
    port map (
      A0 => sig000008b6,
      A1 => sig000008b6,
      A2 => sig000008b6,
      A3 => sig000008b6,
      CE => ce,
      CLK => clk,
      D => sig00000e9a,
      Q => sig00000f79,
      Q15 => NLW_blk0000131a_Q15_UNCONNECTED
    );
  blk0000131b : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => sig00000f79,
      Q => sig00000e7e
    );
  blk0000131c : SRLC16E
    generic map(
      INIT => X"0000"
    )
    port map (
      A0 => sig000008b6,
      A1 => sig000008b6,
      A2 => sig000008b6,
      A3 => sig000008b6,
      CE => ce,
      CLK => clk,
      D => sig00000e99,
      Q => sig00000f7a,
      Q15 => NLW_blk0000131c_Q15_UNCONNECTED
    );
  blk0000131d : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => sig00000f7a,
      Q => sig00000e7d
    );
  blk0000131e : SRLC16E
    generic map(
      INIT => X"0000"
    )
    port map (
      A0 => sig000008b6,
      A1 => sig000008b6,
      A2 => sig000008b6,
      A3 => sig000008b6,
      CE => ce,
      CLK => clk,
      D => sig00000e98,
      Q => sig00000f7b,
      Q15 => NLW_blk0000131e_Q15_UNCONNECTED
    );
  blk0000131f : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => sig00000f7b,
      Q => sig00000e7c
    );
  blk00001320 : SRLC16E
    generic map(
      INIT => X"0000"
    )
    port map (
      A0 => sig000008b6,
      A1 => sig000008b6,
      A2 => sig000008b6,
      A3 => sig000008b6,
      CE => ce,
      CLK => clk,
      D => sig00000e97,
      Q => sig00000f7c,
      Q15 => NLW_blk00001320_Q15_UNCONNECTED
    );
  blk00001321 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => sig00000f7c,
      Q => sig00000e7b
    );
  blk00001322 : SRLC16E
    generic map(
      INIT => X"0000"
    )
    port map (
      A0 => sig000008b6,
      A1 => sig000008b6,
      A2 => sig000008b6,
      A3 => sig000008b6,
      CE => ce,
      CLK => clk,
      D => sig00000e96,
      Q => sig00000f7d,
      Q15 => NLW_blk00001322_Q15_UNCONNECTED
    );
  blk00001323 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => sig00000f7d,
      Q => sig00000e7a
    );
  blk00001324 : SRLC16E
    generic map(
      INIT => X"0000"
    )
    port map (
      A0 => sig000008b6,
      A1 => sig000008b6,
      A2 => sig000008b6,
      A3 => sig000008b6,
      CE => ce,
      CLK => clk,
      D => sig00000e95,
      Q => sig00000f7e,
      Q15 => NLW_blk00001324_Q15_UNCONNECTED
    );
  blk00001325 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => sig00000f7e,
      Q => sig00000e79
    );
  blk00001326 : SRLC16E
    generic map(
      INIT => X"0000"
    )
    port map (
      A0 => sig000008b6,
      A1 => sig000008b6,
      A2 => sig000008b6,
      A3 => sig000008b6,
      CE => ce,
      CLK => clk,
      D => sig00000e94,
      Q => sig00000f7f,
      Q15 => NLW_blk00001326_Q15_UNCONNECTED
    );
  blk00001327 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => sig00000f7f,
      Q => sig00000e78
    );
  blk00001328 : SRLC16E
    generic map(
      INIT => X"0000"
    )
    port map (
      A0 => sig000008b6,
      A1 => sig000008b6,
      A2 => sig000008b6,
      A3 => sig000008b6,
      CE => ce,
      CLK => clk,
      D => sig00000e93,
      Q => sig00000f80,
      Q15 => NLW_blk00001328_Q15_UNCONNECTED
    );
  blk00001329 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => sig00000f80,
      Q => sig00000e77
    );
  blk0000132a : SRLC16E
    generic map(
      INIT => X"0000"
    )
    port map (
      A0 => sig000008b6,
      A1 => sig000008b6,
      A2 => sig000008b6,
      A3 => sig000008b6,
      CE => ce,
      CLK => clk,
      D => sig000000c2,
      Q => sig00000f81,
      Q15 => NLW_blk0000132a_Q15_UNCONNECTED
    );
  blk0000132b : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => sig00000f81,
      Q => sig00000092
    );
  blk0000132c : SRLC16E
    generic map(
      INIT => X"0000"
    )
    port map (
      A0 => sig000008b6,
      A1 => sig000008b6,
      A2 => sig000008b6,
      A3 => sig000008b6,
      CE => ce,
      CLK => clk,
      D => sig000000c1,
      Q => sig00000f82,
      Q15 => NLW_blk0000132c_Q15_UNCONNECTED
    );
  blk0000132d : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => sig00000f82,
      Q => sig00000091
    );
  blk0000132e : SRLC16E
    generic map(
      INIT => X"0000"
    )
    port map (
      A0 => sig000008b6,
      A1 => sig000008b6,
      A2 => sig000008b6,
      A3 => sig000008b6,
      CE => ce,
      CLK => clk,
      D => sig000000c0,
      Q => sig00000f83,
      Q15 => NLW_blk0000132e_Q15_UNCONNECTED
    );
  blk0000132f : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => sig00000f83,
      Q => sig00000090
    );
  blk00001330 : SRLC16E
    generic map(
      INIT => X"0000"
    )
    port map (
      A0 => sig000008b6,
      A1 => sig000008b6,
      A2 => sig000008b6,
      A3 => sig000008b6,
      CE => ce,
      CLK => clk,
      D => sig000000bf,
      Q => sig00000f84,
      Q15 => NLW_blk00001330_Q15_UNCONNECTED
    );
  blk00001331 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => sig00000f84,
      Q => sig0000008f
    );
  blk00001332 : SRLC16E
    generic map(
      INIT => X"0000"
    )
    port map (
      A0 => sig000008b6,
      A1 => sig000008b6,
      A2 => sig000008b6,
      A3 => sig000008b6,
      CE => ce,
      CLK => clk,
      D => sig000000be,
      Q => sig00000f85,
      Q15 => NLW_blk00001332_Q15_UNCONNECTED
    );
  blk00001333 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => sig00000f85,
      Q => sig0000008e
    );
  blk00001334 : SRLC16E
    generic map(
      INIT => X"0000"
    )
    port map (
      A0 => sig000008b6,
      A1 => sig000008b6,
      A2 => sig000008b6,
      A3 => sig000008b6,
      CE => ce,
      CLK => clk,
      D => sig000000bd,
      Q => sig00000f86,
      Q15 => NLW_blk00001334_Q15_UNCONNECTED
    );
  blk00001335 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => sig00000f86,
      Q => sig0000008d
    );
  blk00001336 : SRLC16E
    generic map(
      INIT => X"0000"
    )
    port map (
      A0 => sig000008b6,
      A1 => sig000008b6,
      A2 => sig000008b6,
      A3 => sig000008b6,
      CE => ce,
      CLK => clk,
      D => sig000000bc,
      Q => sig00000f87,
      Q15 => NLW_blk00001336_Q15_UNCONNECTED
    );
  blk00001337 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => sig00000f87,
      Q => sig0000008c
    );
  blk00001338 : SRLC16E
    generic map(
      INIT => X"0000"
    )
    port map (
      A0 => sig000008b6,
      A1 => sig000008b6,
      A2 => sig000008b6,
      A3 => sig000008b6,
      CE => ce,
      CLK => clk,
      D => sig000000bb,
      Q => sig00000f88,
      Q15 => NLW_blk00001338_Q15_UNCONNECTED
    );
  blk00001339 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => sig00000f88,
      Q => sig0000008b
    );
  blk0000133a : SRLC16E
    generic map(
      INIT => X"0000"
    )
    port map (
      A0 => sig000008b6,
      A1 => sig000008b6,
      A2 => sig000008b6,
      A3 => sig000008b6,
      CE => ce,
      CLK => clk,
      D => sig000000ba,
      Q => sig00000f89,
      Q15 => NLW_blk0000133a_Q15_UNCONNECTED
    );
  blk0000133b : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => sig00000f89,
      Q => sig0000008a
    );
  blk0000133c : SRLC16E
    generic map(
      INIT => X"0000"
    )
    port map (
      A0 => sig000008b6,
      A1 => sig000008b6,
      A2 => sig000008b6,
      A3 => sig000008b6,
      CE => ce,
      CLK => clk,
      D => sig000000b9,
      Q => sig00000f8a,
      Q15 => NLW_blk0000133c_Q15_UNCONNECTED
    );
  blk0000133d : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => sig00000f8a,
      Q => sig00000089
    );
  blk0000133e : SRLC16E
    generic map(
      INIT => X"0000"
    )
    port map (
      A0 => sig000008b6,
      A1 => sig000008b6,
      A2 => sig000008b6,
      A3 => sig000008b6,
      CE => ce,
      CLK => clk,
      D => sig000000b8,
      Q => sig00000f8b,
      Q15 => NLW_blk0000133e_Q15_UNCONNECTED
    );
  blk0000133f : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => sig00000f8b,
      Q => sig00000088
    );
  blk00001340 : SRLC16E
    generic map(
      INIT => X"0000"
    )
    port map (
      A0 => sig000008b6,
      A1 => sig000008b6,
      A2 => sig000008b6,
      A3 => sig000008b6,
      CE => ce,
      CLK => clk,
      D => sig000000b7,
      Q => sig00000f8c,
      Q15 => NLW_blk00001340_Q15_UNCONNECTED
    );
  blk00001341 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => sig00000f8c,
      Q => sig00000087
    );
  blk00001342 : SRLC16E
    generic map(
      INIT => X"0000"
    )
    port map (
      A0 => sig000008b6,
      A1 => sig000008b6,
      A2 => sig000008b6,
      A3 => sig000008b6,
      CE => ce,
      CLK => clk,
      D => sig000000b6,
      Q => sig00000f8d,
      Q15 => NLW_blk00001342_Q15_UNCONNECTED
    );
  blk00001343 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => sig00000f8d,
      Q => sig00000086
    );
  blk00001344 : SRLC16E
    generic map(
      INIT => X"0000"
    )
    port map (
      A0 => sig000008b6,
      A1 => sig000008b6,
      A2 => sig000008b6,
      A3 => sig000008b6,
      CE => ce,
      CLK => clk,
      D => sig000000b5,
      Q => sig00000f8e,
      Q15 => NLW_blk00001344_Q15_UNCONNECTED
    );
  blk00001345 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => sig00000f8e,
      Q => sig00000085
    );
  blk00001346 : SRLC16E
    generic map(
      INIT => X"0000"
    )
    port map (
      A0 => sig000008b6,
      A1 => sig000008b6,
      A2 => sig000008b6,
      A3 => sig000008b6,
      CE => ce,
      CLK => clk,
      D => sig000000b4,
      Q => sig00000f8f,
      Q15 => NLW_blk00001346_Q15_UNCONNECTED
    );
  blk00001347 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => sig00000f8f,
      Q => sig00000084
    );
  blk00001348 : SRLC16E
    generic map(
      INIT => X"0000"
    )
    port map (
      A0 => sig000008b6,
      A1 => sig000008b6,
      A2 => sig000008b6,
      A3 => sig000008b6,
      CE => ce,
      CLK => clk,
      D => sig000000b3,
      Q => sig00000f90,
      Q15 => NLW_blk00001348_Q15_UNCONNECTED
    );
  blk00001349 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => sig00000f90,
      Q => sig00000083
    );
  blk0000134a : SRLC16E
    generic map(
      INIT => X"0000"
    )
    port map (
      A0 => sig000008b6,
      A1 => sig000008b6,
      A2 => sig000008b6,
      A3 => sig000008b6,
      CE => ce,
      CLK => clk,
      D => sig000000b2,
      Q => sig00000f91,
      Q15 => NLW_blk0000134a_Q15_UNCONNECTED
    );
  blk0000134b : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => sig00000f91,
      Q => sig00000082
    );
  blk0000134c : SRLC16E
    generic map(
      INIT => X"0000"
    )
    port map (
      A0 => sig000008b6,
      A1 => sig000008b6,
      A2 => sig000008b6,
      A3 => sig000008b6,
      CE => ce,
      CLK => clk,
      D => sig000000b1,
      Q => sig00000f92,
      Q15 => NLW_blk0000134c_Q15_UNCONNECTED
    );
  blk0000134d : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => sig00000f92,
      Q => sig00000081
    );
  blk0000134e : SRLC16E
    generic map(
      INIT => X"0000"
    )
    port map (
      A0 => sig000008b6,
      A1 => sig000008b6,
      A2 => sig000008b6,
      A3 => sig000008b6,
      CE => ce,
      CLK => clk,
      D => sig000000b0,
      Q => sig00000f93,
      Q15 => NLW_blk0000134e_Q15_UNCONNECTED
    );
  blk0000134f : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => sig00000f93,
      Q => sig00000080
    );
  blk00001350 : SRLC16E
    generic map(
      INIT => X"0000"
    )
    port map (
      A0 => sig000008b6,
      A1 => sig000008b6,
      A2 => sig000008b6,
      A3 => sig000008b6,
      CE => ce,
      CLK => clk,
      D => sig000000af,
      Q => sig00000f94,
      Q15 => NLW_blk00001350_Q15_UNCONNECTED
    );
  blk00001351 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => sig00000f94,
      Q => sig0000007f
    );
  blk00001352 : SRLC16E
    generic map(
      INIT => X"0000"
    )
    port map (
      A0 => sig000008b6,
      A1 => sig000008b6,
      A2 => sig000008b6,
      A3 => sig000008b6,
      CE => ce,
      CLK => clk,
      D => sig000000ae,
      Q => sig00000f95,
      Q15 => NLW_blk00001352_Q15_UNCONNECTED
    );
  blk00001353 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => sig00000f95,
      Q => sig0000007e
    );
  blk00001354 : SRLC16E
    generic map(
      INIT => X"0000"
    )
    port map (
      A0 => sig000008b6,
      A1 => sig000008b6,
      A2 => sig000008b6,
      A3 => sig000008b6,
      CE => ce,
      CLK => clk,
      D => sig000000ad,
      Q => sig00000f96,
      Q15 => NLW_blk00001354_Q15_UNCONNECTED
    );
  blk00001355 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => sig00000f96,
      Q => sig0000007d
    );
  blk00001356 : SRLC16E
    generic map(
      INIT => X"0000"
    )
    port map (
      A0 => sig000008b6,
      A1 => sig000008b6,
      A2 => sig000008b6,
      A3 => sig000008b6,
      CE => ce,
      CLK => clk,
      D => sig000000ac,
      Q => sig00000f97,
      Q15 => NLW_blk00001356_Q15_UNCONNECTED
    );
  blk00001357 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => sig00000f97,
      Q => sig0000007c
    );
  blk00001358 : SRLC16E
    generic map(
      INIT => X"0000"
    )
    port map (
      A0 => sig000008b6,
      A1 => sig000008b6,
      A2 => sig000008b6,
      A3 => sig000008b6,
      CE => ce,
      CLK => clk,
      D => sig000000ab,
      Q => sig00000f98,
      Q15 => NLW_blk00001358_Q15_UNCONNECTED
    );
  blk00001359 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => sig00000f98,
      Q => sig0000007b
    );
  blk00000065_blk00000066_blk00000080 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000065_blk00000066_sig00000fdb,
      Q => sig00000140
    );
  blk00000065_blk00000066_blk0000007f : SRLC16E
    generic map(
      INIT => X"0000"
    )
    port map (
      A0 => blk00000065_blk00000066_sig00000fcf,
      A1 => blk00000065_blk00000066_sig00000fce,
      A2 => blk00000065_blk00000066_sig00000fce,
      A3 => blk00000065_blk00000066_sig00000fce,
      CE => ce,
      CLK => clk,
      D => xn_re(10),
      Q => blk00000065_blk00000066_sig00000fdb,
      Q15 => NLW_blk00000065_blk00000066_blk0000007f_Q15_UNCONNECTED
    );
  blk00000065_blk00000066_blk0000007e : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000065_blk00000066_sig00000fda,
      Q => sig0000013f
    );
  blk00000065_blk00000066_blk0000007d : SRLC16E
    generic map(
      INIT => X"0000"
    )
    port map (
      A0 => blk00000065_blk00000066_sig00000fcf,
      A1 => blk00000065_blk00000066_sig00000fce,
      A2 => blk00000065_blk00000066_sig00000fce,
      A3 => blk00000065_blk00000066_sig00000fce,
      CE => ce,
      CLK => clk,
      D => xn_re(9),
      Q => blk00000065_blk00000066_sig00000fda,
      Q15 => NLW_blk00000065_blk00000066_blk0000007d_Q15_UNCONNECTED
    );
  blk00000065_blk00000066_blk0000007c : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000065_blk00000066_sig00000fd9,
      Q => sig00000141
    );
  blk00000065_blk00000066_blk0000007b : SRLC16E
    generic map(
      INIT => X"0000"
    )
    port map (
      A0 => blk00000065_blk00000066_sig00000fcf,
      A1 => blk00000065_blk00000066_sig00000fce,
      A2 => blk00000065_blk00000066_sig00000fce,
      A3 => blk00000065_blk00000066_sig00000fce,
      CE => ce,
      CLK => clk,
      D => xn_re(11),
      Q => blk00000065_blk00000066_sig00000fd9,
      Q15 => NLW_blk00000065_blk00000066_blk0000007b_Q15_UNCONNECTED
    );
  blk00000065_blk00000066_blk0000007a : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000065_blk00000066_sig00000fd8,
      Q => sig0000013d
    );
  blk00000065_blk00000066_blk00000079 : SRLC16E
    generic map(
      INIT => X"0000"
    )
    port map (
      A0 => blk00000065_blk00000066_sig00000fcf,
      A1 => blk00000065_blk00000066_sig00000fce,
      A2 => blk00000065_blk00000066_sig00000fce,
      A3 => blk00000065_blk00000066_sig00000fce,
      CE => ce,
      CLK => clk,
      D => xn_re(7),
      Q => blk00000065_blk00000066_sig00000fd8,
      Q15 => NLW_blk00000065_blk00000066_blk00000079_Q15_UNCONNECTED
    );
  blk00000065_blk00000066_blk00000078 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000065_blk00000066_sig00000fd7,
      Q => sig0000013c
    );
  blk00000065_blk00000066_blk00000077 : SRLC16E
    generic map(
      INIT => X"0000"
    )
    port map (
      A0 => blk00000065_blk00000066_sig00000fcf,
      A1 => blk00000065_blk00000066_sig00000fce,
      A2 => blk00000065_blk00000066_sig00000fce,
      A3 => blk00000065_blk00000066_sig00000fce,
      CE => ce,
      CLK => clk,
      D => xn_re(6),
      Q => blk00000065_blk00000066_sig00000fd7,
      Q15 => NLW_blk00000065_blk00000066_blk00000077_Q15_UNCONNECTED
    );
  blk00000065_blk00000066_blk00000076 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000065_blk00000066_sig00000fd6,
      Q => sig0000013e
    );
  blk00000065_blk00000066_blk00000075 : SRLC16E
    generic map(
      INIT => X"0000"
    )
    port map (
      A0 => blk00000065_blk00000066_sig00000fcf,
      A1 => blk00000065_blk00000066_sig00000fce,
      A2 => blk00000065_blk00000066_sig00000fce,
      A3 => blk00000065_blk00000066_sig00000fce,
      CE => ce,
      CLK => clk,
      D => xn_re(8),
      Q => blk00000065_blk00000066_sig00000fd6,
      Q15 => NLW_blk00000065_blk00000066_blk00000075_Q15_UNCONNECTED
    );
  blk00000065_blk00000066_blk00000074 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000065_blk00000066_sig00000fd5,
      Q => sig0000013a
    );
  blk00000065_blk00000066_blk00000073 : SRLC16E
    generic map(
      INIT => X"0000"
    )
    port map (
      A0 => blk00000065_blk00000066_sig00000fcf,
      A1 => blk00000065_blk00000066_sig00000fce,
      A2 => blk00000065_blk00000066_sig00000fce,
      A3 => blk00000065_blk00000066_sig00000fce,
      CE => ce,
      CLK => clk,
      D => xn_re(4),
      Q => blk00000065_blk00000066_sig00000fd5,
      Q15 => NLW_blk00000065_blk00000066_blk00000073_Q15_UNCONNECTED
    );
  blk00000065_blk00000066_blk00000072 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000065_blk00000066_sig00000fd4,
      Q => sig00000139
    );
  blk00000065_blk00000066_blk00000071 : SRLC16E
    generic map(
      INIT => X"0000"
    )
    port map (
      A0 => blk00000065_blk00000066_sig00000fcf,
      A1 => blk00000065_blk00000066_sig00000fce,
      A2 => blk00000065_blk00000066_sig00000fce,
      A3 => blk00000065_blk00000066_sig00000fce,
      CE => ce,
      CLK => clk,
      D => xn_re(3),
      Q => blk00000065_blk00000066_sig00000fd4,
      Q15 => NLW_blk00000065_blk00000066_blk00000071_Q15_UNCONNECTED
    );
  blk00000065_blk00000066_blk00000070 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000065_blk00000066_sig00000fd3,
      Q => sig0000013b
    );
  blk00000065_blk00000066_blk0000006f : SRLC16E
    generic map(
      INIT => X"0000"
    )
    port map (
      A0 => blk00000065_blk00000066_sig00000fcf,
      A1 => blk00000065_blk00000066_sig00000fce,
      A2 => blk00000065_blk00000066_sig00000fce,
      A3 => blk00000065_blk00000066_sig00000fce,
      CE => ce,
      CLK => clk,
      D => xn_re(5),
      Q => blk00000065_blk00000066_sig00000fd3,
      Q15 => NLW_blk00000065_blk00000066_blk0000006f_Q15_UNCONNECTED
    );
  blk00000065_blk00000066_blk0000006e : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000065_blk00000066_sig00000fd2,
      Q => sig00000137
    );
  blk00000065_blk00000066_blk0000006d : SRLC16E
    generic map(
      INIT => X"0000"
    )
    port map (
      A0 => blk00000065_blk00000066_sig00000fcf,
      A1 => blk00000065_blk00000066_sig00000fce,
      A2 => blk00000065_blk00000066_sig00000fce,
      A3 => blk00000065_blk00000066_sig00000fce,
      CE => ce,
      CLK => clk,
      D => xn_re(1),
      Q => blk00000065_blk00000066_sig00000fd2,
      Q15 => NLW_blk00000065_blk00000066_blk0000006d_Q15_UNCONNECTED
    );
  blk00000065_blk00000066_blk0000006c : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000065_blk00000066_sig00000fd1,
      Q => sig00000136
    );
  blk00000065_blk00000066_blk0000006b : SRLC16E
    generic map(
      INIT => X"0000"
    )
    port map (
      A0 => blk00000065_blk00000066_sig00000fcf,
      A1 => blk00000065_blk00000066_sig00000fce,
      A2 => blk00000065_blk00000066_sig00000fce,
      A3 => blk00000065_blk00000066_sig00000fce,
      CE => ce,
      CLK => clk,
      D => xn_re(0),
      Q => blk00000065_blk00000066_sig00000fd1,
      Q15 => NLW_blk00000065_blk00000066_blk0000006b_Q15_UNCONNECTED
    );
  blk00000065_blk00000066_blk0000006a : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000065_blk00000066_sig00000fd0,
      Q => sig00000138
    );
  blk00000065_blk00000066_blk00000069 : SRLC16E
    generic map(
      INIT => X"0000"
    )
    port map (
      A0 => blk00000065_blk00000066_sig00000fcf,
      A1 => blk00000065_blk00000066_sig00000fce,
      A2 => blk00000065_blk00000066_sig00000fce,
      A3 => blk00000065_blk00000066_sig00000fce,
      CE => ce,
      CLK => clk,
      D => xn_re(2),
      Q => blk00000065_blk00000066_sig00000fd0,
      Q15 => NLW_blk00000065_blk00000066_blk00000069_Q15_UNCONNECTED
    );
  blk00000065_blk00000066_blk00000068 : VCC
    port map (
      P => blk00000065_blk00000066_sig00000fcf
    );
  blk00000065_blk00000066_blk00000067 : GND
    port map (
      G => blk00000065_blk00000066_sig00000fce
    );
  blk00000081_blk00000082_blk0000009c : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000081_blk00000082_sig0000101e,
      Q => sig00000134
    );
  blk00000081_blk00000082_blk0000009b : SRLC16E
    generic map(
      INIT => X"0000"
    )
    port map (
      A0 => blk00000081_blk00000082_sig00001012,
      A1 => blk00000081_blk00000082_sig00001011,
      A2 => blk00000081_blk00000082_sig00001011,
      A3 => blk00000081_blk00000082_sig00001011,
      CE => ce,
      CLK => clk,
      D => xn_im(10),
      Q => blk00000081_blk00000082_sig0000101e,
      Q15 => NLW_blk00000081_blk00000082_blk0000009b_Q15_UNCONNECTED
    );
  blk00000081_blk00000082_blk0000009a : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000081_blk00000082_sig0000101d,
      Q => sig00000133
    );
  blk00000081_blk00000082_blk00000099 : SRLC16E
    generic map(
      INIT => X"0000"
    )
    port map (
      A0 => blk00000081_blk00000082_sig00001012,
      A1 => blk00000081_blk00000082_sig00001011,
      A2 => blk00000081_blk00000082_sig00001011,
      A3 => blk00000081_blk00000082_sig00001011,
      CE => ce,
      CLK => clk,
      D => xn_im(9),
      Q => blk00000081_blk00000082_sig0000101d,
      Q15 => NLW_blk00000081_blk00000082_blk00000099_Q15_UNCONNECTED
    );
  blk00000081_blk00000082_blk00000098 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000081_blk00000082_sig0000101c,
      Q => sig00000135
    );
  blk00000081_blk00000082_blk00000097 : SRLC16E
    generic map(
      INIT => X"0000"
    )
    port map (
      A0 => blk00000081_blk00000082_sig00001012,
      A1 => blk00000081_blk00000082_sig00001011,
      A2 => blk00000081_blk00000082_sig00001011,
      A3 => blk00000081_blk00000082_sig00001011,
      CE => ce,
      CLK => clk,
      D => xn_im(11),
      Q => blk00000081_blk00000082_sig0000101c,
      Q15 => NLW_blk00000081_blk00000082_blk00000097_Q15_UNCONNECTED
    );
  blk00000081_blk00000082_blk00000096 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000081_blk00000082_sig0000101b,
      Q => sig00000131
    );
  blk00000081_blk00000082_blk00000095 : SRLC16E
    generic map(
      INIT => X"0000"
    )
    port map (
      A0 => blk00000081_blk00000082_sig00001012,
      A1 => blk00000081_blk00000082_sig00001011,
      A2 => blk00000081_blk00000082_sig00001011,
      A3 => blk00000081_blk00000082_sig00001011,
      CE => ce,
      CLK => clk,
      D => xn_im(7),
      Q => blk00000081_blk00000082_sig0000101b,
      Q15 => NLW_blk00000081_blk00000082_blk00000095_Q15_UNCONNECTED
    );
  blk00000081_blk00000082_blk00000094 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000081_blk00000082_sig0000101a,
      Q => sig00000130
    );
  blk00000081_blk00000082_blk00000093 : SRLC16E
    generic map(
      INIT => X"0000"
    )
    port map (
      A0 => blk00000081_blk00000082_sig00001012,
      A1 => blk00000081_blk00000082_sig00001011,
      A2 => blk00000081_blk00000082_sig00001011,
      A3 => blk00000081_blk00000082_sig00001011,
      CE => ce,
      CLK => clk,
      D => xn_im(6),
      Q => blk00000081_blk00000082_sig0000101a,
      Q15 => NLW_blk00000081_blk00000082_blk00000093_Q15_UNCONNECTED
    );
  blk00000081_blk00000082_blk00000092 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000081_blk00000082_sig00001019,
      Q => sig00000132
    );
  blk00000081_blk00000082_blk00000091 : SRLC16E
    generic map(
      INIT => X"0000"
    )
    port map (
      A0 => blk00000081_blk00000082_sig00001012,
      A1 => blk00000081_blk00000082_sig00001011,
      A2 => blk00000081_blk00000082_sig00001011,
      A3 => blk00000081_blk00000082_sig00001011,
      CE => ce,
      CLK => clk,
      D => xn_im(8),
      Q => blk00000081_blk00000082_sig00001019,
      Q15 => NLW_blk00000081_blk00000082_blk00000091_Q15_UNCONNECTED
    );
  blk00000081_blk00000082_blk00000090 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000081_blk00000082_sig00001018,
      Q => sig0000012e
    );
  blk00000081_blk00000082_blk0000008f : SRLC16E
    generic map(
      INIT => X"0000"
    )
    port map (
      A0 => blk00000081_blk00000082_sig00001012,
      A1 => blk00000081_blk00000082_sig00001011,
      A2 => blk00000081_blk00000082_sig00001011,
      A3 => blk00000081_blk00000082_sig00001011,
      CE => ce,
      CLK => clk,
      D => xn_im(4),
      Q => blk00000081_blk00000082_sig00001018,
      Q15 => NLW_blk00000081_blk00000082_blk0000008f_Q15_UNCONNECTED
    );
  blk00000081_blk00000082_blk0000008e : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000081_blk00000082_sig00001017,
      Q => sig0000012d
    );
  blk00000081_blk00000082_blk0000008d : SRLC16E
    generic map(
      INIT => X"0000"
    )
    port map (
      A0 => blk00000081_blk00000082_sig00001012,
      A1 => blk00000081_blk00000082_sig00001011,
      A2 => blk00000081_blk00000082_sig00001011,
      A3 => blk00000081_blk00000082_sig00001011,
      CE => ce,
      CLK => clk,
      D => xn_im(3),
      Q => blk00000081_blk00000082_sig00001017,
      Q15 => NLW_blk00000081_blk00000082_blk0000008d_Q15_UNCONNECTED
    );
  blk00000081_blk00000082_blk0000008c : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000081_blk00000082_sig00001016,
      Q => sig0000012f
    );
  blk00000081_blk00000082_blk0000008b : SRLC16E
    generic map(
      INIT => X"0000"
    )
    port map (
      A0 => blk00000081_blk00000082_sig00001012,
      A1 => blk00000081_blk00000082_sig00001011,
      A2 => blk00000081_blk00000082_sig00001011,
      A3 => blk00000081_blk00000082_sig00001011,
      CE => ce,
      CLK => clk,
      D => xn_im(5),
      Q => blk00000081_blk00000082_sig00001016,
      Q15 => NLW_blk00000081_blk00000082_blk0000008b_Q15_UNCONNECTED
    );
  blk00000081_blk00000082_blk0000008a : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000081_blk00000082_sig00001015,
      Q => sig0000012b
    );
  blk00000081_blk00000082_blk00000089 : SRLC16E
    generic map(
      INIT => X"0000"
    )
    port map (
      A0 => blk00000081_blk00000082_sig00001012,
      A1 => blk00000081_blk00000082_sig00001011,
      A2 => blk00000081_blk00000082_sig00001011,
      A3 => blk00000081_blk00000082_sig00001011,
      CE => ce,
      CLK => clk,
      D => xn_im(1),
      Q => blk00000081_blk00000082_sig00001015,
      Q15 => NLW_blk00000081_blk00000082_blk00000089_Q15_UNCONNECTED
    );
  blk00000081_blk00000082_blk00000088 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000081_blk00000082_sig00001014,
      Q => sig0000012a
    );
  blk00000081_blk00000082_blk00000087 : SRLC16E
    generic map(
      INIT => X"0000"
    )
    port map (
      A0 => blk00000081_blk00000082_sig00001012,
      A1 => blk00000081_blk00000082_sig00001011,
      A2 => blk00000081_blk00000082_sig00001011,
      A3 => blk00000081_blk00000082_sig00001011,
      CE => ce,
      CLK => clk,
      D => xn_im(0),
      Q => blk00000081_blk00000082_sig00001014,
      Q15 => NLW_blk00000081_blk00000082_blk00000087_Q15_UNCONNECTED
    );
  blk00000081_blk00000082_blk00000086 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000081_blk00000082_sig00001013,
      Q => sig0000012c
    );
  blk00000081_blk00000082_blk00000085 : SRLC16E
    generic map(
      INIT => X"0000"
    )
    port map (
      A0 => blk00000081_blk00000082_sig00001012,
      A1 => blk00000081_blk00000082_sig00001011,
      A2 => blk00000081_blk00000082_sig00001011,
      A3 => blk00000081_blk00000082_sig00001011,
      CE => ce,
      CLK => clk,
      D => xn_im(2),
      Q => blk00000081_blk00000082_sig00001013,
      Q15 => NLW_blk00000081_blk00000082_blk00000085_Q15_UNCONNECTED
    );
  blk00000081_blk00000082_blk00000084 : VCC
    port map (
      P => blk00000081_blk00000082_sig00001012
    );
  blk00000081_blk00000082_blk00000083 : GND
    port map (
      G => blk00000081_blk00000082_sig00001011
    );
  blk000000ed_blk00000103 : LUT1
    generic map(
      INIT => X"2"
    )
    port map (
      I0 => sig00000165,
      O => blk000000ed_sig0000103e
    );
  blk000000ed_blk00000102 : LUT1
    generic map(
      INIT => X"2"
    )
    port map (
      I0 => sig00000164,
      O => blk000000ed_sig0000103d
    );
  blk000000ed_blk00000101 : LUT1
    generic map(
      INIT => X"2"
    )
    port map (
      I0 => sig00000163,
      O => blk000000ed_sig0000103c
    );
  blk000000ed_blk00000100 : LUT1
    generic map(
      INIT => X"2"
    )
    port map (
      I0 => sig00000162,
      O => blk000000ed_sig0000103b
    );
  blk000000ed_blk000000ff : LUT1
    generic map(
      INIT => X"2"
    )
    port map (
      I0 => sig00000161,
      O => blk000000ed_sig0000103a
    );
  blk000000ed_blk000000fe : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => sig00000186,
      D => blk000000ed_sig00001038,
      R => sig000008b6,
      Q => NlwRenamedSig_OI_xn_index(0)
    );
  blk000000ed_blk000000fd : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => sig00000186,
      D => blk000000ed_sig00001033,
      R => sig000008b6,
      Q => NlwRenamedSig_OI_xn_index(1)
    );
  blk000000ed_blk000000fc : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => sig00000186,
      D => blk000000ed_sig00001032,
      R => sig000008b6,
      Q => NlwRenamedSig_OI_xn_index(2)
    );
  blk000000ed_blk000000fb : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => sig00000186,
      D => blk000000ed_sig00001031,
      R => sig000008b6,
      Q => NlwRenamedSig_OI_xn_index(3)
    );
  blk000000ed_blk000000fa : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => sig00000186,
      D => blk000000ed_sig00001030,
      R => sig000008b6,
      Q => NlwRenamedSig_OI_xn_index(4)
    );
  blk000000ed_blk000000f9 : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => sig00000186,
      D => blk000000ed_sig0000102f,
      R => sig000008b6,
      Q => NlwRenamedSig_OI_xn_index(5)
    );
  blk000000ed_blk000000f8 : MUXCY
    port map (
      CI => sig00000167,
      DI => sig00000165,
      S => blk000000ed_sig0000103e,
      O => blk000000ed_sig00001039
    );
  blk000000ed_blk000000f7 : XORCY
    port map (
      CI => sig00000167,
      LI => blk000000ed_sig0000103e,
      O => blk000000ed_sig00001038
    );
  blk000000ed_blk000000f6 : MUXCY
    port map (
      CI => blk000000ed_sig00001039,
      DI => sig00000164,
      S => blk000000ed_sig0000103d,
      O => blk000000ed_sig00001037
    );
  blk000000ed_blk000000f5 : MUXCY
    port map (
      CI => blk000000ed_sig00001037,
      DI => sig00000163,
      S => blk000000ed_sig0000103c,
      O => blk000000ed_sig00001036
    );
  blk000000ed_blk000000f4 : MUXCY
    port map (
      CI => blk000000ed_sig00001036,
      DI => sig00000162,
      S => blk000000ed_sig0000103b,
      O => blk000000ed_sig00001035
    );
  blk000000ed_blk000000f3 : MUXCY
    port map (
      CI => blk000000ed_sig00001035,
      DI => sig00000161,
      S => blk000000ed_sig0000103a,
      O => blk000000ed_sig00001034
    );
  blk000000ed_blk000000f2 : XORCY
    port map (
      CI => blk000000ed_sig00001039,
      LI => blk000000ed_sig0000103d,
      O => blk000000ed_sig00001033
    );
  blk000000ed_blk000000f1 : XORCY
    port map (
      CI => blk000000ed_sig00001037,
      LI => blk000000ed_sig0000103c,
      O => blk000000ed_sig00001032
    );
  blk000000ed_blk000000f0 : XORCY
    port map (
      CI => blk000000ed_sig00001036,
      LI => blk000000ed_sig0000103b,
      O => blk000000ed_sig00001031
    );
  blk000000ed_blk000000ef : XORCY
    port map (
      CI => blk000000ed_sig00001035,
      LI => blk000000ed_sig0000103a,
      O => blk000000ed_sig00001030
    );
  blk000000ed_blk000000ee : XORCY
    port map (
      CI => blk000000ed_sig00001034,
      LI => sig00000160,
      O => blk000000ed_sig0000102f
    );
  blk00000104_blk0000011a : LUT1
    generic map(
      INIT => X"2"
    )
    port map (
      I0 => sig0000001b,
      O => blk00000104_sig0000105e
    );
  blk00000104_blk00000119 : LUT1
    generic map(
      INIT => X"2"
    )
    port map (
      I0 => sig0000001c,
      O => blk00000104_sig0000105d
    );
  blk00000104_blk00000118 : LUT1
    generic map(
      INIT => X"2"
    )
    port map (
      I0 => sig0000001d,
      O => blk00000104_sig0000105c
    );
  blk00000104_blk00000117 : LUT1
    generic map(
      INIT => X"2"
    )
    port map (
      I0 => sig0000001e,
      O => blk00000104_sig0000105b
    );
  blk00000104_blk00000116 : LUT1
    generic map(
      INIT => X"2"
    )
    port map (
      I0 => sig0000001f,
      O => blk00000104_sig0000105a
    );
  blk00000104_blk00000115 : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => sig00000017,
      D => blk00000104_sig00001058,
      R => sig000008b6,
      Q => sig0000011b
    );
  blk00000104_blk00000114 : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => sig00000017,
      D => blk00000104_sig00001053,
      R => sig000008b6,
      Q => sig0000011a
    );
  blk00000104_blk00000113 : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => sig00000017,
      D => blk00000104_sig00001052,
      R => sig000008b6,
      Q => sig00000119
    );
  blk00000104_blk00000112 : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => sig00000017,
      D => blk00000104_sig00001051,
      R => sig000008b6,
      Q => sig00000118
    );
  blk00000104_blk00000111 : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => sig00000017,
      D => blk00000104_sig00001050,
      R => sig000008b6,
      Q => sig00000117
    );
  blk00000104_blk00000110 : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => sig00000017,
      D => blk00000104_sig0000104f,
      R => sig000008b6,
      Q => sig00000116
    );
  blk00000104_blk0000010f : MUXCY
    port map (
      CI => sig00000019,
      DI => sig0000001b,
      S => blk00000104_sig0000105e,
      O => blk00000104_sig00001059
    );
  blk00000104_blk0000010e : XORCY
    port map (
      CI => sig00000019,
      LI => blk00000104_sig0000105e,
      O => blk00000104_sig00001058
    );
  blk00000104_blk0000010d : MUXCY
    port map (
      CI => blk00000104_sig00001059,
      DI => sig0000001c,
      S => blk00000104_sig0000105d,
      O => blk00000104_sig00001057
    );
  blk00000104_blk0000010c : MUXCY
    port map (
      CI => blk00000104_sig00001057,
      DI => sig0000001d,
      S => blk00000104_sig0000105c,
      O => blk00000104_sig00001056
    );
  blk00000104_blk0000010b : MUXCY
    port map (
      CI => blk00000104_sig00001056,
      DI => sig0000001e,
      S => blk00000104_sig0000105b,
      O => blk00000104_sig00001055
    );
  blk00000104_blk0000010a : MUXCY
    port map (
      CI => blk00000104_sig00001055,
      DI => sig0000001f,
      S => blk00000104_sig0000105a,
      O => blk00000104_sig00001054
    );
  blk00000104_blk00000109 : XORCY
    port map (
      CI => blk00000104_sig00001059,
      LI => blk00000104_sig0000105d,
      O => blk00000104_sig00001053
    );
  blk00000104_blk00000108 : XORCY
    port map (
      CI => blk00000104_sig00001057,
      LI => blk00000104_sig0000105c,
      O => blk00000104_sig00001052
    );
  blk00000104_blk00000107 : XORCY
    port map (
      CI => blk00000104_sig00001056,
      LI => blk00000104_sig0000105b,
      O => blk00000104_sig00001051
    );
  blk00000104_blk00000106 : XORCY
    port map (
      CI => blk00000104_sig00001055,
      LI => blk00000104_sig0000105a,
      O => blk00000104_sig00001050
    );
  blk00000104_blk00000105 : XORCY
    port map (
      CI => blk00000104_sig00001054,
      LI => sig00000020,
      O => blk00000104_sig0000104f
    );
  blk0000011b_blk00000131 : LUT1
    generic map(
      INIT => X"2"
    )
    port map (
      I0 => sig000001bf,
      O => blk0000011b_sig0000107e
    );
  blk0000011b_blk00000130 : LUT1
    generic map(
      INIT => X"2"
    )
    port map (
      I0 => sig000001c0,
      O => blk0000011b_sig0000107d
    );
  blk0000011b_blk0000012f : LUT1
    generic map(
      INIT => X"2"
    )
    port map (
      I0 => sig000001c1,
      O => blk0000011b_sig0000107c
    );
  blk0000011b_blk0000012e : LUT1
    generic map(
      INIT => X"2"
    )
    port map (
      I0 => sig000001c2,
      O => blk0000011b_sig0000107b
    );
  blk0000011b_blk0000012d : LUT1
    generic map(
      INIT => X"2"
    )
    port map (
      I0 => sig000001c3,
      O => blk0000011b_sig0000107a
    );
  blk0000011b_blk0000012c : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => sig00000185,
      D => blk0000011b_sig00001078,
      R => sig000008b6,
      Q => sig00000192
    );
  blk0000011b_blk0000012b : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => sig00000185,
      D => blk0000011b_sig00001073,
      R => sig000008b6,
      Q => sig00000193
    );
  blk0000011b_blk0000012a : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => sig00000185,
      D => blk0000011b_sig00001072,
      R => sig000008b6,
      Q => sig00000194
    );
  blk0000011b_blk00000129 : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => sig00000185,
      D => blk0000011b_sig00001071,
      R => sig000008b6,
      Q => sig00000195
    );
  blk0000011b_blk00000128 : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => sig00000185,
      D => blk0000011b_sig00001070,
      R => sig000008b6,
      Q => sig00000196
    );
  blk0000011b_blk00000127 : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => sig00000185,
      D => blk0000011b_sig0000106f,
      R => sig000008b6,
      Q => sig00000197
    );
  blk0000011b_blk00000126 : MUXCY
    port map (
      CI => sig000001b9,
      DI => sig000001bf,
      S => blk0000011b_sig0000107e,
      O => blk0000011b_sig00001079
    );
  blk0000011b_blk00000125 : XORCY
    port map (
      CI => sig000001b9,
      LI => blk0000011b_sig0000107e,
      O => blk0000011b_sig00001078
    );
  blk0000011b_blk00000124 : MUXCY
    port map (
      CI => blk0000011b_sig00001079,
      DI => sig000001c0,
      S => blk0000011b_sig0000107d,
      O => blk0000011b_sig00001077
    );
  blk0000011b_blk00000123 : MUXCY
    port map (
      CI => blk0000011b_sig00001077,
      DI => sig000001c1,
      S => blk0000011b_sig0000107c,
      O => blk0000011b_sig00001076
    );
  blk0000011b_blk00000122 : MUXCY
    port map (
      CI => blk0000011b_sig00001076,
      DI => sig000001c2,
      S => blk0000011b_sig0000107b,
      O => blk0000011b_sig00001075
    );
  blk0000011b_blk00000121 : MUXCY
    port map (
      CI => blk0000011b_sig00001075,
      DI => sig000001c3,
      S => blk0000011b_sig0000107a,
      O => blk0000011b_sig00001074
    );
  blk0000011b_blk00000120 : XORCY
    port map (
      CI => blk0000011b_sig00001079,
      LI => blk0000011b_sig0000107d,
      O => blk0000011b_sig00001073
    );
  blk0000011b_blk0000011f : XORCY
    port map (
      CI => blk0000011b_sig00001077,
      LI => blk0000011b_sig0000107c,
      O => blk0000011b_sig00001072
    );
  blk0000011b_blk0000011e : XORCY
    port map (
      CI => blk0000011b_sig00001076,
      LI => blk0000011b_sig0000107b,
      O => blk0000011b_sig00001071
    );
  blk0000011b_blk0000011d : XORCY
    port map (
      CI => blk0000011b_sig00001075,
      LI => blk0000011b_sig0000107a,
      O => blk0000011b_sig00001070
    );
  blk0000011b_blk0000011c : XORCY
    port map (
      CI => blk0000011b_sig00001074,
      LI => sig000001c4,
      O => blk0000011b_sig0000106f
    );
  blk0000014b_blk00000161 : LUT1
    generic map(
      INIT => X"2"
    )
    port map (
      I0 => sig000001e0,
      O => blk0000014b_sig0000109e
    );
  blk0000014b_blk00000160 : LUT1
    generic map(
      INIT => X"2"
    )
    port map (
      I0 => sig000001e1,
      O => blk0000014b_sig0000109d
    );
  blk0000014b_blk0000015f : LUT1
    generic map(
      INIT => X"2"
    )
    port map (
      I0 => sig000001e2,
      O => blk0000014b_sig0000109c
    );
  blk0000014b_blk0000015e : LUT1
    generic map(
      INIT => X"2"
    )
    port map (
      I0 => sig000001e3,
      O => blk0000014b_sig0000109b
    );
  blk0000014b_blk0000015d : LUT1
    generic map(
      INIT => X"2"
    )
    port map (
      I0 => sig000001e4,
      O => blk0000014b_sig0000109a
    );
  blk0000014b_blk0000015c : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => sig00000013,
      D => blk0000014b_sig00001098,
      R => sig000008b6,
      Q => sig000000a4
    );
  blk0000014b_blk0000015b : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => sig00000013,
      D => blk0000014b_sig00001093,
      R => sig000008b6,
      Q => sig000000a5
    );
  blk0000014b_blk0000015a : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => sig00000013,
      D => blk0000014b_sig00001092,
      R => sig000008b6,
      Q => sig000000a6
    );
  blk0000014b_blk00000159 : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => sig00000013,
      D => blk0000014b_sig00001091,
      R => sig000008b6,
      Q => sig000000a7
    );
  blk0000014b_blk00000158 : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => sig00000013,
      D => blk0000014b_sig00001090,
      R => sig000008b6,
      Q => sig000000a8
    );
  blk0000014b_blk00000157 : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => sig00000013,
      D => blk0000014b_sig0000108f,
      R => sig000008b6,
      Q => sig000000a9
    );
  blk0000014b_blk00000156 : MUXCY
    port map (
      CI => sig000001da,
      DI => sig000001e0,
      S => blk0000014b_sig0000109e,
      O => blk0000014b_sig00001099
    );
  blk0000014b_blk00000155 : XORCY
    port map (
      CI => sig000001da,
      LI => blk0000014b_sig0000109e,
      O => blk0000014b_sig00001098
    );
  blk0000014b_blk00000154 : MUXCY
    port map (
      CI => blk0000014b_sig00001099,
      DI => sig000001e1,
      S => blk0000014b_sig0000109d,
      O => blk0000014b_sig00001097
    );
  blk0000014b_blk00000153 : MUXCY
    port map (
      CI => blk0000014b_sig00001097,
      DI => sig000001e2,
      S => blk0000014b_sig0000109c,
      O => blk0000014b_sig00001096
    );
  blk0000014b_blk00000152 : MUXCY
    port map (
      CI => blk0000014b_sig00001096,
      DI => sig000001e3,
      S => blk0000014b_sig0000109b,
      O => blk0000014b_sig00001095
    );
  blk0000014b_blk00000151 : MUXCY
    port map (
      CI => blk0000014b_sig00001095,
      DI => sig000001e4,
      S => blk0000014b_sig0000109a,
      O => blk0000014b_sig00001094
    );
  blk0000014b_blk00000150 : XORCY
    port map (
      CI => blk0000014b_sig00001099,
      LI => blk0000014b_sig0000109d,
      O => blk0000014b_sig00001093
    );
  blk0000014b_blk0000014f : XORCY
    port map (
      CI => blk0000014b_sig00001097,
      LI => blk0000014b_sig0000109c,
      O => blk0000014b_sig00001092
    );
  blk0000014b_blk0000014e : XORCY
    port map (
      CI => blk0000014b_sig00001096,
      LI => blk0000014b_sig0000109b,
      O => blk0000014b_sig00001091
    );
  blk0000014b_blk0000014d : XORCY
    port map (
      CI => blk0000014b_sig00001095,
      LI => blk0000014b_sig0000109a,
      O => blk0000014b_sig00001090
    );
  blk0000014b_blk0000014c : XORCY
    port map (
      CI => blk0000014b_sig00001094,
      LI => sig000001e5,
      O => blk0000014b_sig0000108f
    );
  blk0000017b_blk0000017c_blk00000180 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk0000017b_blk0000017c_sig000010b0,
      Q => sig00000190
    );
  blk0000017b_blk0000017c_blk0000017f : SRLC16E
    generic map(
      INIT => X"0000"
    )
    port map (
      A0 => blk0000017b_blk0000017c_sig000010af,
      A1 => blk0000017b_blk0000017c_sig000010ae,
      A2 => blk0000017b_blk0000017c_sig000010ae,
      A3 => blk0000017b_blk0000017c_sig000010ae,
      CE => ce,
      CLK => clk,
      D => sig0000018b,
      Q => blk0000017b_blk0000017c_sig000010b0,
      Q15 => NLW_blk0000017b_blk0000017c_blk0000017f_Q15_UNCONNECTED
    );
  blk0000017b_blk0000017c_blk0000017e : VCC
    port map (
      P => blk0000017b_blk0000017c_sig000010af
    );
  blk0000017b_blk0000017c_blk0000017d : GND
    port map (
      G => blk0000017b_blk0000017c_sig000010ae
    );
  blk00000181_blk00000182_blk00000186 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000181_blk00000182_sig000010c2,
      Q => sig00000005
    );
  blk00000181_blk00000182_blk00000185 : SRLC16E
    generic map(
      INIT => X"0000"
    )
    port map (
      A0 => blk00000181_blk00000182_sig000010c1,
      A1 => blk00000181_blk00000182_sig000010c0,
      A2 => blk00000181_blk00000182_sig000010c0,
      A3 => blk00000181_blk00000182_sig000010c0,
      CE => ce,
      CLK => clk,
      D => sig00000048,
      Q => blk00000181_blk00000182_sig000010c2,
      Q15 => NLW_blk00000181_blk00000182_blk00000185_Q15_UNCONNECTED
    );
  blk00000181_blk00000182_blk00000184 : VCC
    port map (
      P => blk00000181_blk00000182_sig000010c1
    );
  blk00000181_blk00000182_blk00000183 : GND
    port map (
      G => blk00000181_blk00000182_sig000010c0
    );
  blk00000187_blk00000188_blk0000018c : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000187_blk00000188_sig000010d4,
      Q => sig00000003
    );
  blk00000187_blk00000188_blk0000018b : SRLC16E
    generic map(
      INIT => X"0000"
    )
    port map (
      A0 => blk00000187_blk00000188_sig000010d3,
      A1 => blk00000187_blk00000188_sig000010d2,
      A2 => blk00000187_blk00000188_sig000010d2,
      A3 => blk00000187_blk00000188_sig000010d2,
      CE => ce,
      CLK => clk,
      D => sig00000114,
      Q => blk00000187_blk00000188_sig000010d4,
      Q15 => NLW_blk00000187_blk00000188_blk0000018b_Q15_UNCONNECTED
    );
  blk00000187_blk00000188_blk0000018a : VCC
    port map (
      P => blk00000187_blk00000188_sig000010d3
    );
  blk00000187_blk00000188_blk00000189 : GND
    port map (
      G => blk00000187_blk00000188_sig000010d2
    );
  blk0000018d_blk0000018e_blk00000192 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk0000018d_blk0000018e_sig000010ea,
      Q => sig00000113
    );
  blk0000018d_blk0000018e_blk00000191 : SRLC16E
    generic map(
      INIT => X"0000"
    )
    port map (
      A0 => blk0000018d_blk0000018e_sig000010e9,
      A1 => blk0000018d_blk0000018e_sig000010e8,
      A2 => blk0000018d_blk0000018e_sig000010e8,
      A3 => blk0000018d_blk0000018e_sig000010e8,
      CE => ce,
      CLK => clk,
      D => NlwRenamedSig_OI_xn_index(5),
      Q => blk0000018d_blk0000018e_sig000010ea,
      Q15 => NLW_blk0000018d_blk0000018e_blk00000191_Q15_UNCONNECTED
    );
  blk0000018d_blk0000018e_blk00000190 : VCC
    port map (
      P => blk0000018d_blk0000018e_sig000010e9
    );
  blk0000018d_blk0000018e_blk0000018f : GND
    port map (
      G => blk0000018d_blk0000018e_sig000010e8
    );
  blk00000193_blk00000194_blk0000019a : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000193_blk00000194_sig00001103,
      Q => sig00000250
    );
  blk00000193_blk00000194_blk00000199 : SRLC16E
    generic map(
      INIT => X"0000"
    )
    port map (
      A0 => blk00000193_blk00000194_sig00001101,
      A1 => blk00000193_blk00000194_sig00001100,
      A2 => blk00000193_blk00000194_sig00001100,
      A3 => blk00000193_blk00000194_sig00001100,
      CE => ce,
      CLK => clk,
      D => sig00000288,
      Q => blk00000193_blk00000194_sig00001103,
      Q15 => NLW_blk00000193_blk00000194_blk00000199_Q15_UNCONNECTED
    );
  blk00000193_blk00000194_blk00000198 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000193_blk00000194_sig00001102,
      Q => sig0000024f
    );
  blk00000193_blk00000194_blk00000197 : SRLC16E
    generic map(
      INIT => X"0000"
    )
    port map (
      A0 => blk00000193_blk00000194_sig00001101,
      A1 => blk00000193_blk00000194_sig00001100,
      A2 => blk00000193_blk00000194_sig00001100,
      A3 => blk00000193_blk00000194_sig00001100,
      CE => ce,
      CLK => clk,
      D => sig00000287,
      Q => blk00000193_blk00000194_sig00001102,
      Q15 => NLW_blk00000193_blk00000194_blk00000197_Q15_UNCONNECTED
    );
  blk00000193_blk00000194_blk00000196 : VCC
    port map (
      P => blk00000193_blk00000194_sig00001101
    );
  blk00000193_blk00000194_blk00000195 : GND
    port map (
      G => blk00000193_blk00000194_sig00001100
    );
  blk000001aa_blk000001c0 : LUT1
    generic map(
      INIT => X"2"
    )
    port map (
      I0 => sig00000297,
      O => blk000001aa_sig00001123
    );
  blk000001aa_blk000001bf : LUT1
    generic map(
      INIT => X"2"
    )
    port map (
      I0 => sig00000296,
      O => blk000001aa_sig00001122
    );
  blk000001aa_blk000001be : LUT1
    generic map(
      INIT => X"2"
    )
    port map (
      I0 => sig00000295,
      O => blk000001aa_sig00001121
    );
  blk000001aa_blk000001bd : LUT1
    generic map(
      INIT => X"2"
    )
    port map (
      I0 => sig00000294,
      O => blk000001aa_sig00001120
    );
  blk000001aa_blk000001bc : LUT1
    generic map(
      INIT => X"2"
    )
    port map (
      I0 => sig00000293,
      O => blk000001aa_sig0000111f
    );
  blk000001aa_blk000001bb : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => sig0000029e,
      D => blk000001aa_sig0000111d,
      R => sig000008b6,
      Q => sig00000283
    );
  blk000001aa_blk000001ba : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => sig0000029e,
      D => blk000001aa_sig00001118,
      R => sig000008b6,
      Q => sig00000284
    );
  blk000001aa_blk000001b9 : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => sig0000029e,
      D => blk000001aa_sig00001117,
      R => sig000008b6,
      Q => sig00000285
    );
  blk000001aa_blk000001b8 : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => sig0000029e,
      D => blk000001aa_sig00001116,
      R => sig000008b6,
      Q => sig00000286
    );
  blk000001aa_blk000001b7 : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => sig0000029e,
      D => blk000001aa_sig00001115,
      R => sig000008b6,
      Q => sig00000287
    );
  blk000001aa_blk000001b6 : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => sig0000029e,
      D => blk000001aa_sig00001114,
      R => sig000008b6,
      Q => sig00000288
    );
  blk000001aa_blk000001b5 : MUXCY
    port map (
      CI => sig00000299,
      DI => sig00000297,
      S => blk000001aa_sig00001123,
      O => blk000001aa_sig0000111e
    );
  blk000001aa_blk000001b4 : XORCY
    port map (
      CI => sig00000299,
      LI => blk000001aa_sig00001123,
      O => blk000001aa_sig0000111d
    );
  blk000001aa_blk000001b3 : MUXCY
    port map (
      CI => blk000001aa_sig0000111e,
      DI => sig00000296,
      S => blk000001aa_sig00001122,
      O => blk000001aa_sig0000111c
    );
  blk000001aa_blk000001b2 : MUXCY
    port map (
      CI => blk000001aa_sig0000111c,
      DI => sig00000295,
      S => blk000001aa_sig00001121,
      O => blk000001aa_sig0000111b
    );
  blk000001aa_blk000001b1 : MUXCY
    port map (
      CI => blk000001aa_sig0000111b,
      DI => sig00000294,
      S => blk000001aa_sig00001120,
      O => blk000001aa_sig0000111a
    );
  blk000001aa_blk000001b0 : MUXCY
    port map (
      CI => blk000001aa_sig0000111a,
      DI => sig00000293,
      S => blk000001aa_sig0000111f,
      O => blk000001aa_sig00001119
    );
  blk000001aa_blk000001af : XORCY
    port map (
      CI => blk000001aa_sig0000111e,
      LI => blk000001aa_sig00001122,
      O => blk000001aa_sig00001118
    );
  blk000001aa_blk000001ae : XORCY
    port map (
      CI => blk000001aa_sig0000111c,
      LI => blk000001aa_sig00001121,
      O => blk000001aa_sig00001117
    );
  blk000001aa_blk000001ad : XORCY
    port map (
      CI => blk000001aa_sig0000111b,
      LI => blk000001aa_sig00001120,
      O => blk000001aa_sig00001116
    );
  blk000001aa_blk000001ac : XORCY
    port map (
      CI => blk000001aa_sig0000111a,
      LI => blk000001aa_sig0000111f,
      O => blk000001aa_sig00001115
    );
  blk000001aa_blk000001ab : XORCY
    port map (
      CI => blk000001aa_sig00001119,
      LI => sig00000292,
      O => blk000001aa_sig00001114
    );
  blk000001d2_blk000001e8 : LUT1
    generic map(
      INIT => X"2"
    )
    port map (
      I0 => sig000002af,
      O => blk000001d2_sig00001143
    );
  blk000001d2_blk000001e7 : LUT1
    generic map(
      INIT => X"2"
    )
    port map (
      I0 => sig000002ae,
      O => blk000001d2_sig00001142
    );
  blk000001d2_blk000001e6 : LUT1
    generic map(
      INIT => X"2"
    )
    port map (
      I0 => sig000002ad,
      O => blk000001d2_sig00001141
    );
  blk000001d2_blk000001e5 : LUT1
    generic map(
      INIT => X"2"
    )
    port map (
      I0 => sig000002ac,
      O => blk000001d2_sig00001140
    );
  blk000001d2_blk000001e4 : LUT1
    generic map(
      INIT => X"2"
    )
    port map (
      I0 => sig000002ab,
      O => blk000001d2_sig0000113f
    );
  blk000001d2_blk000001e3 : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => sig000002b6,
      D => blk000001d2_sig0000113d,
      R => sig000008b6,
      Q => sig0000027c
    );
  blk000001d2_blk000001e2 : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => sig000002b6,
      D => blk000001d2_sig00001138,
      R => sig000008b6,
      Q => sig0000027d
    );
  blk000001d2_blk000001e1 : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => sig000002b6,
      D => blk000001d2_sig00001137,
      R => sig000008b6,
      Q => sig0000027e
    );
  blk000001d2_blk000001e0 : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => sig000002b6,
      D => blk000001d2_sig00001136,
      R => sig000008b6,
      Q => sig0000027f
    );
  blk000001d2_blk000001df : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => sig000002b6,
      D => blk000001d2_sig00001135,
      R => sig000008b6,
      Q => sig00000280
    );
  blk000001d2_blk000001de : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => sig000002b6,
      D => blk000001d2_sig00001134,
      R => sig000008b6,
      Q => sig00000281
    );
  blk000001d2_blk000001dd : MUXCY
    port map (
      CI => sig000002b1,
      DI => sig000002af,
      S => blk000001d2_sig00001143,
      O => blk000001d2_sig0000113e
    );
  blk000001d2_blk000001dc : XORCY
    port map (
      CI => sig000002b1,
      LI => blk000001d2_sig00001143,
      O => blk000001d2_sig0000113d
    );
  blk000001d2_blk000001db : MUXCY
    port map (
      CI => blk000001d2_sig0000113e,
      DI => sig000002ae,
      S => blk000001d2_sig00001142,
      O => blk000001d2_sig0000113c
    );
  blk000001d2_blk000001da : MUXCY
    port map (
      CI => blk000001d2_sig0000113c,
      DI => sig000002ad,
      S => blk000001d2_sig00001141,
      O => blk000001d2_sig0000113b
    );
  blk000001d2_blk000001d9 : MUXCY
    port map (
      CI => blk000001d2_sig0000113b,
      DI => sig000002ac,
      S => blk000001d2_sig00001140,
      O => blk000001d2_sig0000113a
    );
  blk000001d2_blk000001d8 : MUXCY
    port map (
      CI => blk000001d2_sig0000113a,
      DI => sig000002ab,
      S => blk000001d2_sig0000113f,
      O => blk000001d2_sig00001139
    );
  blk000001d2_blk000001d7 : XORCY
    port map (
      CI => blk000001d2_sig0000113e,
      LI => blk000001d2_sig00001142,
      O => blk000001d2_sig00001138
    );
  blk000001d2_blk000001d6 : XORCY
    port map (
      CI => blk000001d2_sig0000113c,
      LI => blk000001d2_sig00001141,
      O => blk000001d2_sig00001137
    );
  blk000001d2_blk000001d5 : XORCY
    port map (
      CI => blk000001d2_sig0000113b,
      LI => blk000001d2_sig00001140,
      O => blk000001d2_sig00001136
    );
  blk000001d2_blk000001d4 : XORCY
    port map (
      CI => blk000001d2_sig0000113a,
      LI => blk000001d2_sig0000113f,
      O => blk000001d2_sig00001135
    );
  blk000001d2_blk000001d3 : XORCY
    port map (
      CI => blk000001d2_sig00001139,
      LI => sig000002aa,
      O => blk000001d2_sig00001134
    );
  blk000001fa_blk000001fb_blk000001ff : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk000001fa_blk000001fb_sig00001155,
      Q => sig0000030c
    );
  blk000001fa_blk000001fb_blk000001fe : SRLC16E
    generic map(
      INIT => X"0000"
    )
    port map (
      A0 => blk000001fa_blk000001fb_sig00001154,
      A1 => blk000001fa_blk000001fb_sig00001153,
      A2 => blk000001fa_blk000001fb_sig00001153,
      A3 => blk000001fa_blk000001fb_sig00001153,
      CE => ce,
      CLK => clk,
      D => sig00000113,
      Q => blk000001fa_blk000001fb_sig00001155,
      Q15 => NLW_blk000001fa_blk000001fb_blk000001fe_Q15_UNCONNECTED
    );
  blk000001fa_blk000001fb_blk000001fd : VCC
    port map (
      P => blk000001fa_blk000001fb_sig00001154
    );
  blk000001fa_blk000001fb_blk000001fc : GND
    port map (
      G => blk000001fa_blk000001fb_sig00001153
    );
  blk00000200_blk00000201_blk0000021b : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000200_blk00000201_sig00001198,
      Q => sig00000317
    );
  blk00000200_blk00000201_blk0000021a : SRLC16E
    generic map(
      INIT => X"0000"
    )
    port map (
      A0 => blk00000200_blk00000201_sig0000118c,
      A1 => blk00000200_blk00000201_sig0000118b,
      A2 => blk00000200_blk00000201_sig0000118b,
      A3 => blk00000200_blk00000201_sig0000118b,
      CE => ce,
      CLK => clk,
      D => sig00000134,
      Q => blk00000200_blk00000201_sig00001198,
      Q15 => NLW_blk00000200_blk00000201_blk0000021a_Q15_UNCONNECTED
    );
  blk00000200_blk00000201_blk00000219 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000200_blk00000201_sig00001197,
      Q => sig00000316
    );
  blk00000200_blk00000201_blk00000218 : SRLC16E
    generic map(
      INIT => X"0000"
    )
    port map (
      A0 => blk00000200_blk00000201_sig0000118c,
      A1 => blk00000200_blk00000201_sig0000118b,
      A2 => blk00000200_blk00000201_sig0000118b,
      A3 => blk00000200_blk00000201_sig0000118b,
      CE => ce,
      CLK => clk,
      D => sig00000133,
      Q => blk00000200_blk00000201_sig00001197,
      Q15 => NLW_blk00000200_blk00000201_blk00000218_Q15_UNCONNECTED
    );
  blk00000200_blk00000201_blk00000217 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000200_blk00000201_sig00001196,
      Q => sig00000318
    );
  blk00000200_blk00000201_blk00000216 : SRLC16E
    generic map(
      INIT => X"0000"
    )
    port map (
      A0 => blk00000200_blk00000201_sig0000118c,
      A1 => blk00000200_blk00000201_sig0000118b,
      A2 => blk00000200_blk00000201_sig0000118b,
      A3 => blk00000200_blk00000201_sig0000118b,
      CE => ce,
      CLK => clk,
      D => sig00000135,
      Q => blk00000200_blk00000201_sig00001196,
      Q15 => NLW_blk00000200_blk00000201_blk00000216_Q15_UNCONNECTED
    );
  blk00000200_blk00000201_blk00000215 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000200_blk00000201_sig00001195,
      Q => sig00000314
    );
  blk00000200_blk00000201_blk00000214 : SRLC16E
    generic map(
      INIT => X"0000"
    )
    port map (
      A0 => blk00000200_blk00000201_sig0000118c,
      A1 => blk00000200_blk00000201_sig0000118b,
      A2 => blk00000200_blk00000201_sig0000118b,
      A3 => blk00000200_blk00000201_sig0000118b,
      CE => ce,
      CLK => clk,
      D => sig00000131,
      Q => blk00000200_blk00000201_sig00001195,
      Q15 => NLW_blk00000200_blk00000201_blk00000214_Q15_UNCONNECTED
    );
  blk00000200_blk00000201_blk00000213 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000200_blk00000201_sig00001194,
      Q => sig00000313
    );
  blk00000200_blk00000201_blk00000212 : SRLC16E
    generic map(
      INIT => X"0000"
    )
    port map (
      A0 => blk00000200_blk00000201_sig0000118c,
      A1 => blk00000200_blk00000201_sig0000118b,
      A2 => blk00000200_blk00000201_sig0000118b,
      A3 => blk00000200_blk00000201_sig0000118b,
      CE => ce,
      CLK => clk,
      D => sig00000130,
      Q => blk00000200_blk00000201_sig00001194,
      Q15 => NLW_blk00000200_blk00000201_blk00000212_Q15_UNCONNECTED
    );
  blk00000200_blk00000201_blk00000211 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000200_blk00000201_sig00001193,
      Q => sig00000315
    );
  blk00000200_blk00000201_blk00000210 : SRLC16E
    generic map(
      INIT => X"0000"
    )
    port map (
      A0 => blk00000200_blk00000201_sig0000118c,
      A1 => blk00000200_blk00000201_sig0000118b,
      A2 => blk00000200_blk00000201_sig0000118b,
      A3 => blk00000200_blk00000201_sig0000118b,
      CE => ce,
      CLK => clk,
      D => sig00000132,
      Q => blk00000200_blk00000201_sig00001193,
      Q15 => NLW_blk00000200_blk00000201_blk00000210_Q15_UNCONNECTED
    );
  blk00000200_blk00000201_blk0000020f : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000200_blk00000201_sig00001192,
      Q => sig00000311
    );
  blk00000200_blk00000201_blk0000020e : SRLC16E
    generic map(
      INIT => X"0000"
    )
    port map (
      A0 => blk00000200_blk00000201_sig0000118c,
      A1 => blk00000200_blk00000201_sig0000118b,
      A2 => blk00000200_blk00000201_sig0000118b,
      A3 => blk00000200_blk00000201_sig0000118b,
      CE => ce,
      CLK => clk,
      D => sig0000012e,
      Q => blk00000200_blk00000201_sig00001192,
      Q15 => NLW_blk00000200_blk00000201_blk0000020e_Q15_UNCONNECTED
    );
  blk00000200_blk00000201_blk0000020d : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000200_blk00000201_sig00001191,
      Q => sig00000310
    );
  blk00000200_blk00000201_blk0000020c : SRLC16E
    generic map(
      INIT => X"0000"
    )
    port map (
      A0 => blk00000200_blk00000201_sig0000118c,
      A1 => blk00000200_blk00000201_sig0000118b,
      A2 => blk00000200_blk00000201_sig0000118b,
      A3 => blk00000200_blk00000201_sig0000118b,
      CE => ce,
      CLK => clk,
      D => sig0000012d,
      Q => blk00000200_blk00000201_sig00001191,
      Q15 => NLW_blk00000200_blk00000201_blk0000020c_Q15_UNCONNECTED
    );
  blk00000200_blk00000201_blk0000020b : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000200_blk00000201_sig00001190,
      Q => sig00000312
    );
  blk00000200_blk00000201_blk0000020a : SRLC16E
    generic map(
      INIT => X"0000"
    )
    port map (
      A0 => blk00000200_blk00000201_sig0000118c,
      A1 => blk00000200_blk00000201_sig0000118b,
      A2 => blk00000200_blk00000201_sig0000118b,
      A3 => blk00000200_blk00000201_sig0000118b,
      CE => ce,
      CLK => clk,
      D => sig0000012f,
      Q => blk00000200_blk00000201_sig00001190,
      Q15 => NLW_blk00000200_blk00000201_blk0000020a_Q15_UNCONNECTED
    );
  blk00000200_blk00000201_blk00000209 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000200_blk00000201_sig0000118f,
      Q => sig0000030e
    );
  blk00000200_blk00000201_blk00000208 : SRLC16E
    generic map(
      INIT => X"0000"
    )
    port map (
      A0 => blk00000200_blk00000201_sig0000118c,
      A1 => blk00000200_blk00000201_sig0000118b,
      A2 => blk00000200_blk00000201_sig0000118b,
      A3 => blk00000200_blk00000201_sig0000118b,
      CE => ce,
      CLK => clk,
      D => sig0000012b,
      Q => blk00000200_blk00000201_sig0000118f,
      Q15 => NLW_blk00000200_blk00000201_blk00000208_Q15_UNCONNECTED
    );
  blk00000200_blk00000201_blk00000207 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000200_blk00000201_sig0000118e,
      Q => sig0000030d
    );
  blk00000200_blk00000201_blk00000206 : SRLC16E
    generic map(
      INIT => X"0000"
    )
    port map (
      A0 => blk00000200_blk00000201_sig0000118c,
      A1 => blk00000200_blk00000201_sig0000118b,
      A2 => blk00000200_blk00000201_sig0000118b,
      A3 => blk00000200_blk00000201_sig0000118b,
      CE => ce,
      CLK => clk,
      D => sig0000012a,
      Q => blk00000200_blk00000201_sig0000118e,
      Q15 => NLW_blk00000200_blk00000201_blk00000206_Q15_UNCONNECTED
    );
  blk00000200_blk00000201_blk00000205 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000200_blk00000201_sig0000118d,
      Q => sig0000030f
    );
  blk00000200_blk00000201_blk00000204 : SRLC16E
    generic map(
      INIT => X"0000"
    )
    port map (
      A0 => blk00000200_blk00000201_sig0000118c,
      A1 => blk00000200_blk00000201_sig0000118b,
      A2 => blk00000200_blk00000201_sig0000118b,
      A3 => blk00000200_blk00000201_sig0000118b,
      CE => ce,
      CLK => clk,
      D => sig0000012c,
      Q => blk00000200_blk00000201_sig0000118d,
      Q15 => NLW_blk00000200_blk00000201_blk00000204_Q15_UNCONNECTED
    );
  blk00000200_blk00000201_blk00000203 : VCC
    port map (
      P => blk00000200_blk00000201_sig0000118c
    );
  blk00000200_blk00000201_blk00000202 : GND
    port map (
      G => blk00000200_blk00000201_sig0000118b
    );
  blk0000021c_blk0000021d_blk00000237 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk0000021c_blk0000021d_sig000011db,
      Q => sig00000323
    );
  blk0000021c_blk0000021d_blk00000236 : SRLC16E
    generic map(
      INIT => X"0000"
    )
    port map (
      A0 => blk0000021c_blk0000021d_sig000011cf,
      A1 => blk0000021c_blk0000021d_sig000011ce,
      A2 => blk0000021c_blk0000021d_sig000011ce,
      A3 => blk0000021c_blk0000021d_sig000011ce,
      CE => ce,
      CLK => clk,
      D => sig00000140,
      Q => blk0000021c_blk0000021d_sig000011db,
      Q15 => NLW_blk0000021c_blk0000021d_blk00000236_Q15_UNCONNECTED
    );
  blk0000021c_blk0000021d_blk00000235 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk0000021c_blk0000021d_sig000011da,
      Q => sig00000322
    );
  blk0000021c_blk0000021d_blk00000234 : SRLC16E
    generic map(
      INIT => X"0000"
    )
    port map (
      A0 => blk0000021c_blk0000021d_sig000011cf,
      A1 => blk0000021c_blk0000021d_sig000011ce,
      A2 => blk0000021c_blk0000021d_sig000011ce,
      A3 => blk0000021c_blk0000021d_sig000011ce,
      CE => ce,
      CLK => clk,
      D => sig0000013f,
      Q => blk0000021c_blk0000021d_sig000011da,
      Q15 => NLW_blk0000021c_blk0000021d_blk00000234_Q15_UNCONNECTED
    );
  blk0000021c_blk0000021d_blk00000233 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk0000021c_blk0000021d_sig000011d9,
      Q => sig00000324
    );
  blk0000021c_blk0000021d_blk00000232 : SRLC16E
    generic map(
      INIT => X"0000"
    )
    port map (
      A0 => blk0000021c_blk0000021d_sig000011cf,
      A1 => blk0000021c_blk0000021d_sig000011ce,
      A2 => blk0000021c_blk0000021d_sig000011ce,
      A3 => blk0000021c_blk0000021d_sig000011ce,
      CE => ce,
      CLK => clk,
      D => sig00000141,
      Q => blk0000021c_blk0000021d_sig000011d9,
      Q15 => NLW_blk0000021c_blk0000021d_blk00000232_Q15_UNCONNECTED
    );
  blk0000021c_blk0000021d_blk00000231 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk0000021c_blk0000021d_sig000011d8,
      Q => sig00000320
    );
  blk0000021c_blk0000021d_blk00000230 : SRLC16E
    generic map(
      INIT => X"0000"
    )
    port map (
      A0 => blk0000021c_blk0000021d_sig000011cf,
      A1 => blk0000021c_blk0000021d_sig000011ce,
      A2 => blk0000021c_blk0000021d_sig000011ce,
      A3 => blk0000021c_blk0000021d_sig000011ce,
      CE => ce,
      CLK => clk,
      D => sig0000013d,
      Q => blk0000021c_blk0000021d_sig000011d8,
      Q15 => NLW_blk0000021c_blk0000021d_blk00000230_Q15_UNCONNECTED
    );
  blk0000021c_blk0000021d_blk0000022f : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk0000021c_blk0000021d_sig000011d7,
      Q => sig0000031f
    );
  blk0000021c_blk0000021d_blk0000022e : SRLC16E
    generic map(
      INIT => X"0000"
    )
    port map (
      A0 => blk0000021c_blk0000021d_sig000011cf,
      A1 => blk0000021c_blk0000021d_sig000011ce,
      A2 => blk0000021c_blk0000021d_sig000011ce,
      A3 => blk0000021c_blk0000021d_sig000011ce,
      CE => ce,
      CLK => clk,
      D => sig0000013c,
      Q => blk0000021c_blk0000021d_sig000011d7,
      Q15 => NLW_blk0000021c_blk0000021d_blk0000022e_Q15_UNCONNECTED
    );
  blk0000021c_blk0000021d_blk0000022d : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk0000021c_blk0000021d_sig000011d6,
      Q => sig00000321
    );
  blk0000021c_blk0000021d_blk0000022c : SRLC16E
    generic map(
      INIT => X"0000"
    )
    port map (
      A0 => blk0000021c_blk0000021d_sig000011cf,
      A1 => blk0000021c_blk0000021d_sig000011ce,
      A2 => blk0000021c_blk0000021d_sig000011ce,
      A3 => blk0000021c_blk0000021d_sig000011ce,
      CE => ce,
      CLK => clk,
      D => sig0000013e,
      Q => blk0000021c_blk0000021d_sig000011d6,
      Q15 => NLW_blk0000021c_blk0000021d_blk0000022c_Q15_UNCONNECTED
    );
  blk0000021c_blk0000021d_blk0000022b : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk0000021c_blk0000021d_sig000011d5,
      Q => sig0000031d
    );
  blk0000021c_blk0000021d_blk0000022a : SRLC16E
    generic map(
      INIT => X"0000"
    )
    port map (
      A0 => blk0000021c_blk0000021d_sig000011cf,
      A1 => blk0000021c_blk0000021d_sig000011ce,
      A2 => blk0000021c_blk0000021d_sig000011ce,
      A3 => blk0000021c_blk0000021d_sig000011ce,
      CE => ce,
      CLK => clk,
      D => sig0000013a,
      Q => blk0000021c_blk0000021d_sig000011d5,
      Q15 => NLW_blk0000021c_blk0000021d_blk0000022a_Q15_UNCONNECTED
    );
  blk0000021c_blk0000021d_blk00000229 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk0000021c_blk0000021d_sig000011d4,
      Q => sig0000031c
    );
  blk0000021c_blk0000021d_blk00000228 : SRLC16E
    generic map(
      INIT => X"0000"
    )
    port map (
      A0 => blk0000021c_blk0000021d_sig000011cf,
      A1 => blk0000021c_blk0000021d_sig000011ce,
      A2 => blk0000021c_blk0000021d_sig000011ce,
      A3 => blk0000021c_blk0000021d_sig000011ce,
      CE => ce,
      CLK => clk,
      D => sig00000139,
      Q => blk0000021c_blk0000021d_sig000011d4,
      Q15 => NLW_blk0000021c_blk0000021d_blk00000228_Q15_UNCONNECTED
    );
  blk0000021c_blk0000021d_blk00000227 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk0000021c_blk0000021d_sig000011d3,
      Q => sig0000031e
    );
  blk0000021c_blk0000021d_blk00000226 : SRLC16E
    generic map(
      INIT => X"0000"
    )
    port map (
      A0 => blk0000021c_blk0000021d_sig000011cf,
      A1 => blk0000021c_blk0000021d_sig000011ce,
      A2 => blk0000021c_blk0000021d_sig000011ce,
      A3 => blk0000021c_blk0000021d_sig000011ce,
      CE => ce,
      CLK => clk,
      D => sig0000013b,
      Q => blk0000021c_blk0000021d_sig000011d3,
      Q15 => NLW_blk0000021c_blk0000021d_blk00000226_Q15_UNCONNECTED
    );
  blk0000021c_blk0000021d_blk00000225 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk0000021c_blk0000021d_sig000011d2,
      Q => sig0000031a
    );
  blk0000021c_blk0000021d_blk00000224 : SRLC16E
    generic map(
      INIT => X"0000"
    )
    port map (
      A0 => blk0000021c_blk0000021d_sig000011cf,
      A1 => blk0000021c_blk0000021d_sig000011ce,
      A2 => blk0000021c_blk0000021d_sig000011ce,
      A3 => blk0000021c_blk0000021d_sig000011ce,
      CE => ce,
      CLK => clk,
      D => sig00000137,
      Q => blk0000021c_blk0000021d_sig000011d2,
      Q15 => NLW_blk0000021c_blk0000021d_blk00000224_Q15_UNCONNECTED
    );
  blk0000021c_blk0000021d_blk00000223 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk0000021c_blk0000021d_sig000011d1,
      Q => sig00000319
    );
  blk0000021c_blk0000021d_blk00000222 : SRLC16E
    generic map(
      INIT => X"0000"
    )
    port map (
      A0 => blk0000021c_blk0000021d_sig000011cf,
      A1 => blk0000021c_blk0000021d_sig000011ce,
      A2 => blk0000021c_blk0000021d_sig000011ce,
      A3 => blk0000021c_blk0000021d_sig000011ce,
      CE => ce,
      CLK => clk,
      D => sig00000136,
      Q => blk0000021c_blk0000021d_sig000011d1,
      Q15 => NLW_blk0000021c_blk0000021d_blk00000222_Q15_UNCONNECTED
    );
  blk0000021c_blk0000021d_blk00000221 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk0000021c_blk0000021d_sig000011d0,
      Q => sig0000031b
    );
  blk0000021c_blk0000021d_blk00000220 : SRLC16E
    generic map(
      INIT => X"0000"
    )
    port map (
      A0 => blk0000021c_blk0000021d_sig000011cf,
      A1 => blk0000021c_blk0000021d_sig000011ce,
      A2 => blk0000021c_blk0000021d_sig000011ce,
      A3 => blk0000021c_blk0000021d_sig000011ce,
      CE => ce,
      CLK => clk,
      D => sig00000138,
      Q => blk0000021c_blk0000021d_sig000011d0,
      Q15 => NLW_blk0000021c_blk0000021d_blk00000220_Q15_UNCONNECTED
    );
  blk0000021c_blk0000021d_blk0000021f : VCC
    port map (
      P => blk0000021c_blk0000021d_sig000011cf
    );
  blk0000021c_blk0000021d_blk0000021e : GND
    port map (
      G => blk0000021c_blk0000021d_sig000011ce
    );
  blk00000287_blk00000288_blk000002be : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000287_blk00000288_sig00001263,
      Q => sig000002ef
    );
  blk00000287_blk00000288_blk000002bd : SRLC32E
    generic map(
      INIT => X"00000000"
    )
    port map (
      CLK => clk,
      D => sig00000309,
      CE => ce,
      Q => blk00000287_blk00000288_sig00001263,
      Q31 => NLW_blk00000287_blk00000288_blk000002bd_Q31_UNCONNECTED,
      A(4) => blk00000287_blk00000288_sig00001249,
      A(3) => blk00000287_blk00000288_sig00001249,
      A(2) => blk00000287_blk00000288_sig00001249,
      A(1) => blk00000287_blk00000288_sig00001248,
      A(0) => blk00000287_blk00000288_sig00001248
    );
  blk00000287_blk00000288_blk000002bc : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000287_blk00000288_sig00001262,
      Q => sig000002ee
    );
  blk00000287_blk00000288_blk000002bb : SRLC32E
    generic map(
      INIT => X"00000000"
    )
    port map (
      CLK => clk,
      D => sig00000308,
      CE => ce,
      Q => blk00000287_blk00000288_sig00001262,
      Q31 => NLW_blk00000287_blk00000288_blk000002bb_Q31_UNCONNECTED,
      A(4) => blk00000287_blk00000288_sig00001249,
      A(3) => blk00000287_blk00000288_sig00001249,
      A(2) => blk00000287_blk00000288_sig00001249,
      A(1) => blk00000287_blk00000288_sig00001248,
      A(0) => blk00000287_blk00000288_sig00001248
    );
  blk00000287_blk00000288_blk000002ba : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000287_blk00000288_sig00001261,
      Q => sig000002f0
    );
  blk00000287_blk00000288_blk000002b9 : SRLC32E
    generic map(
      INIT => X"00000000"
    )
    port map (
      CLK => clk,
      D => sig0000030a,
      CE => ce,
      Q => blk00000287_blk00000288_sig00001261,
      Q31 => NLW_blk00000287_blk00000288_blk000002b9_Q31_UNCONNECTED,
      A(4) => blk00000287_blk00000288_sig00001249,
      A(3) => blk00000287_blk00000288_sig00001249,
      A(2) => blk00000287_blk00000288_sig00001249,
      A(1) => blk00000287_blk00000288_sig00001248,
      A(0) => blk00000287_blk00000288_sig00001248
    );
  blk00000287_blk00000288_blk000002b8 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000287_blk00000288_sig00001260,
      Q => sig000002ec
    );
  blk00000287_blk00000288_blk000002b7 : SRLC32E
    generic map(
      INIT => X"00000000"
    )
    port map (
      CLK => clk,
      D => sig00000306,
      CE => ce,
      Q => blk00000287_blk00000288_sig00001260,
      Q31 => NLW_blk00000287_blk00000288_blk000002b7_Q31_UNCONNECTED,
      A(4) => blk00000287_blk00000288_sig00001249,
      A(3) => blk00000287_blk00000288_sig00001249,
      A(2) => blk00000287_blk00000288_sig00001249,
      A(1) => blk00000287_blk00000288_sig00001248,
      A(0) => blk00000287_blk00000288_sig00001248
    );
  blk00000287_blk00000288_blk000002b6 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000287_blk00000288_sig0000125f,
      Q => sig000002eb
    );
  blk00000287_blk00000288_blk000002b5 : SRLC32E
    generic map(
      INIT => X"00000000"
    )
    port map (
      CLK => clk,
      D => sig00000305,
      CE => ce,
      Q => blk00000287_blk00000288_sig0000125f,
      Q31 => NLW_blk00000287_blk00000288_blk000002b5_Q31_UNCONNECTED,
      A(4) => blk00000287_blk00000288_sig00001249,
      A(3) => blk00000287_blk00000288_sig00001249,
      A(2) => blk00000287_blk00000288_sig00001249,
      A(1) => blk00000287_blk00000288_sig00001248,
      A(0) => blk00000287_blk00000288_sig00001248
    );
  blk00000287_blk00000288_blk000002b4 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000287_blk00000288_sig0000125e,
      Q => sig000002ed
    );
  blk00000287_blk00000288_blk000002b3 : SRLC32E
    generic map(
      INIT => X"00000000"
    )
    port map (
      CLK => clk,
      D => sig00000307,
      CE => ce,
      Q => blk00000287_blk00000288_sig0000125e,
      Q31 => NLW_blk00000287_blk00000288_blk000002b3_Q31_UNCONNECTED,
      A(4) => blk00000287_blk00000288_sig00001249,
      A(3) => blk00000287_blk00000288_sig00001249,
      A(2) => blk00000287_blk00000288_sig00001249,
      A(1) => blk00000287_blk00000288_sig00001248,
      A(0) => blk00000287_blk00000288_sig00001248
    );
  blk00000287_blk00000288_blk000002b2 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000287_blk00000288_sig0000125d,
      Q => sig000002e9
    );
  blk00000287_blk00000288_blk000002b1 : SRLC32E
    generic map(
      INIT => X"00000000"
    )
    port map (
      CLK => clk,
      D => sig00000303,
      CE => ce,
      Q => blk00000287_blk00000288_sig0000125d,
      Q31 => NLW_blk00000287_blk00000288_blk000002b1_Q31_UNCONNECTED,
      A(4) => blk00000287_blk00000288_sig00001249,
      A(3) => blk00000287_blk00000288_sig00001249,
      A(2) => blk00000287_blk00000288_sig00001249,
      A(1) => blk00000287_blk00000288_sig00001248,
      A(0) => blk00000287_blk00000288_sig00001248
    );
  blk00000287_blk00000288_blk000002b0 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000287_blk00000288_sig0000125c,
      Q => sig000002e8
    );
  blk00000287_blk00000288_blk000002af : SRLC32E
    generic map(
      INIT => X"00000000"
    )
    port map (
      CLK => clk,
      D => sig00000302,
      CE => ce,
      Q => blk00000287_blk00000288_sig0000125c,
      Q31 => NLW_blk00000287_blk00000288_blk000002af_Q31_UNCONNECTED,
      A(4) => blk00000287_blk00000288_sig00001249,
      A(3) => blk00000287_blk00000288_sig00001249,
      A(2) => blk00000287_blk00000288_sig00001249,
      A(1) => blk00000287_blk00000288_sig00001248,
      A(0) => blk00000287_blk00000288_sig00001248
    );
  blk00000287_blk00000288_blk000002ae : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000287_blk00000288_sig0000125b,
      Q => sig000002ea
    );
  blk00000287_blk00000288_blk000002ad : SRLC32E
    generic map(
      INIT => X"00000000"
    )
    port map (
      CLK => clk,
      D => sig00000304,
      CE => ce,
      Q => blk00000287_blk00000288_sig0000125b,
      Q31 => NLW_blk00000287_blk00000288_blk000002ad_Q31_UNCONNECTED,
      A(4) => blk00000287_blk00000288_sig00001249,
      A(3) => blk00000287_blk00000288_sig00001249,
      A(2) => blk00000287_blk00000288_sig00001249,
      A(1) => blk00000287_blk00000288_sig00001248,
      A(0) => blk00000287_blk00000288_sig00001248
    );
  blk00000287_blk00000288_blk000002ac : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000287_blk00000288_sig0000125a,
      Q => sig000002e7
    );
  blk00000287_blk00000288_blk000002ab : SRLC32E
    generic map(
      INIT => X"00000000"
    )
    port map (
      CLK => clk,
      D => sig00000301,
      CE => ce,
      Q => blk00000287_blk00000288_sig0000125a,
      Q31 => NLW_blk00000287_blk00000288_blk000002ab_Q31_UNCONNECTED,
      A(4) => blk00000287_blk00000288_sig00001249,
      A(3) => blk00000287_blk00000288_sig00001249,
      A(2) => blk00000287_blk00000288_sig00001249,
      A(1) => blk00000287_blk00000288_sig00001248,
      A(0) => blk00000287_blk00000288_sig00001248
    );
  blk00000287_blk00000288_blk000002aa : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000287_blk00000288_sig00001259,
      Q => sig000002e6
    );
  blk00000287_blk00000288_blk000002a9 : SRLC32E
    generic map(
      INIT => X"00000000"
    )
    port map (
      CLK => clk,
      D => sig00000300,
      CE => ce,
      Q => blk00000287_blk00000288_sig00001259,
      Q31 => NLW_blk00000287_blk00000288_blk000002a9_Q31_UNCONNECTED,
      A(4) => blk00000287_blk00000288_sig00001249,
      A(3) => blk00000287_blk00000288_sig00001249,
      A(2) => blk00000287_blk00000288_sig00001249,
      A(1) => blk00000287_blk00000288_sig00001248,
      A(0) => blk00000287_blk00000288_sig00001248
    );
  blk00000287_blk00000288_blk000002a8 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000287_blk00000288_sig00001258,
      Q => sig000002e5
    );
  blk00000287_blk00000288_blk000002a7 : SRLC32E
    generic map(
      INIT => X"00000000"
    )
    port map (
      CLK => clk,
      D => sig000002ff,
      CE => ce,
      Q => blk00000287_blk00000288_sig00001258,
      Q31 => NLW_blk00000287_blk00000288_blk000002a7_Q31_UNCONNECTED,
      A(4) => blk00000287_blk00000288_sig00001249,
      A(3) => blk00000287_blk00000288_sig00001249,
      A(2) => blk00000287_blk00000288_sig00001249,
      A(1) => blk00000287_blk00000288_sig00001248,
      A(0) => blk00000287_blk00000288_sig00001248
    );
  blk00000287_blk00000288_blk000002a6 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000287_blk00000288_sig00001257,
      Q => sig000002e4
    );
  blk00000287_blk00000288_blk000002a5 : SRLC32E
    generic map(
      INIT => X"00000000"
    )
    port map (
      CLK => clk,
      D => sig000002fe,
      CE => ce,
      Q => blk00000287_blk00000288_sig00001257,
      Q31 => NLW_blk00000287_blk00000288_blk000002a5_Q31_UNCONNECTED,
      A(4) => blk00000287_blk00000288_sig00001249,
      A(3) => blk00000287_blk00000288_sig00001249,
      A(2) => blk00000287_blk00000288_sig00001249,
      A(1) => blk00000287_blk00000288_sig00001248,
      A(0) => blk00000287_blk00000288_sig00001248
    );
  blk00000287_blk00000288_blk000002a4 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000287_blk00000288_sig00001256,
      Q => sig000002e2
    );
  blk00000287_blk00000288_blk000002a3 : SRLC32E
    generic map(
      INIT => X"00000000"
    )
    port map (
      CLK => clk,
      D => sig000002fc,
      CE => ce,
      Q => blk00000287_blk00000288_sig00001256,
      Q31 => NLW_blk00000287_blk00000288_blk000002a3_Q31_UNCONNECTED,
      A(4) => blk00000287_blk00000288_sig00001249,
      A(3) => blk00000287_blk00000288_sig00001249,
      A(2) => blk00000287_blk00000288_sig00001249,
      A(1) => blk00000287_blk00000288_sig00001248,
      A(0) => blk00000287_blk00000288_sig00001248
    );
  blk00000287_blk00000288_blk000002a2 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000287_blk00000288_sig00001255,
      Q => sig000002e1
    );
  blk00000287_blk00000288_blk000002a1 : SRLC32E
    generic map(
      INIT => X"00000000"
    )
    port map (
      CLK => clk,
      D => sig000002fb,
      CE => ce,
      Q => blk00000287_blk00000288_sig00001255,
      Q31 => NLW_blk00000287_blk00000288_blk000002a1_Q31_UNCONNECTED,
      A(4) => blk00000287_blk00000288_sig00001249,
      A(3) => blk00000287_blk00000288_sig00001249,
      A(2) => blk00000287_blk00000288_sig00001249,
      A(1) => blk00000287_blk00000288_sig00001248,
      A(0) => blk00000287_blk00000288_sig00001248
    );
  blk00000287_blk00000288_blk000002a0 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000287_blk00000288_sig00001254,
      Q => sig000002e3
    );
  blk00000287_blk00000288_blk0000029f : SRLC32E
    generic map(
      INIT => X"00000000"
    )
    port map (
      CLK => clk,
      D => sig000002fd,
      CE => ce,
      Q => blk00000287_blk00000288_sig00001254,
      Q31 => NLW_blk00000287_blk00000288_blk0000029f_Q31_UNCONNECTED,
      A(4) => blk00000287_blk00000288_sig00001249,
      A(3) => blk00000287_blk00000288_sig00001249,
      A(2) => blk00000287_blk00000288_sig00001249,
      A(1) => blk00000287_blk00000288_sig00001248,
      A(0) => blk00000287_blk00000288_sig00001248
    );
  blk00000287_blk00000288_blk0000029e : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000287_blk00000288_sig00001253,
      Q => sig000002df
    );
  blk00000287_blk00000288_blk0000029d : SRLC32E
    generic map(
      INIT => X"00000000"
    )
    port map (
      CLK => clk,
      D => sig000002f9,
      CE => ce,
      Q => blk00000287_blk00000288_sig00001253,
      Q31 => NLW_blk00000287_blk00000288_blk0000029d_Q31_UNCONNECTED,
      A(4) => blk00000287_blk00000288_sig00001249,
      A(3) => blk00000287_blk00000288_sig00001249,
      A(2) => blk00000287_blk00000288_sig00001249,
      A(1) => blk00000287_blk00000288_sig00001248,
      A(0) => blk00000287_blk00000288_sig00001248
    );
  blk00000287_blk00000288_blk0000029c : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000287_blk00000288_sig00001252,
      Q => sig000002de
    );
  blk00000287_blk00000288_blk0000029b : SRLC32E
    generic map(
      INIT => X"00000000"
    )
    port map (
      CLK => clk,
      D => sig000002f8,
      CE => ce,
      Q => blk00000287_blk00000288_sig00001252,
      Q31 => NLW_blk00000287_blk00000288_blk0000029b_Q31_UNCONNECTED,
      A(4) => blk00000287_blk00000288_sig00001249,
      A(3) => blk00000287_blk00000288_sig00001249,
      A(2) => blk00000287_blk00000288_sig00001249,
      A(1) => blk00000287_blk00000288_sig00001248,
      A(0) => blk00000287_blk00000288_sig00001248
    );
  blk00000287_blk00000288_blk0000029a : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000287_blk00000288_sig00001251,
      Q => sig000002e0
    );
  blk00000287_blk00000288_blk00000299 : SRLC32E
    generic map(
      INIT => X"00000000"
    )
    port map (
      CLK => clk,
      D => sig000002fa,
      CE => ce,
      Q => blk00000287_blk00000288_sig00001251,
      Q31 => NLW_blk00000287_blk00000288_blk00000299_Q31_UNCONNECTED,
      A(4) => blk00000287_blk00000288_sig00001249,
      A(3) => blk00000287_blk00000288_sig00001249,
      A(2) => blk00000287_blk00000288_sig00001249,
      A(1) => blk00000287_blk00000288_sig00001248,
      A(0) => blk00000287_blk00000288_sig00001248
    );
  blk00000287_blk00000288_blk00000298 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000287_blk00000288_sig00001250,
      Q => sig000002dc
    );
  blk00000287_blk00000288_blk00000297 : SRLC32E
    generic map(
      INIT => X"00000000"
    )
    port map (
      CLK => clk,
      D => sig000002f6,
      CE => ce,
      Q => blk00000287_blk00000288_sig00001250,
      Q31 => NLW_blk00000287_blk00000288_blk00000297_Q31_UNCONNECTED,
      A(4) => blk00000287_blk00000288_sig00001249,
      A(3) => blk00000287_blk00000288_sig00001249,
      A(2) => blk00000287_blk00000288_sig00001249,
      A(1) => blk00000287_blk00000288_sig00001248,
      A(0) => blk00000287_blk00000288_sig00001248
    );
  blk00000287_blk00000288_blk00000296 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000287_blk00000288_sig0000124f,
      Q => sig000002db
    );
  blk00000287_blk00000288_blk00000295 : SRLC32E
    generic map(
      INIT => X"00000000"
    )
    port map (
      CLK => clk,
      D => sig000002f5,
      CE => ce,
      Q => blk00000287_blk00000288_sig0000124f,
      Q31 => NLW_blk00000287_blk00000288_blk00000295_Q31_UNCONNECTED,
      A(4) => blk00000287_blk00000288_sig00001249,
      A(3) => blk00000287_blk00000288_sig00001249,
      A(2) => blk00000287_blk00000288_sig00001249,
      A(1) => blk00000287_blk00000288_sig00001248,
      A(0) => blk00000287_blk00000288_sig00001248
    );
  blk00000287_blk00000288_blk00000294 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000287_blk00000288_sig0000124e,
      Q => sig000002dd
    );
  blk00000287_blk00000288_blk00000293 : SRLC32E
    generic map(
      INIT => X"00000000"
    )
    port map (
      CLK => clk,
      D => sig000002f7,
      CE => ce,
      Q => blk00000287_blk00000288_sig0000124e,
      Q31 => NLW_blk00000287_blk00000288_blk00000293_Q31_UNCONNECTED,
      A(4) => blk00000287_blk00000288_sig00001249,
      A(3) => blk00000287_blk00000288_sig00001249,
      A(2) => blk00000287_blk00000288_sig00001249,
      A(1) => blk00000287_blk00000288_sig00001248,
      A(0) => blk00000287_blk00000288_sig00001248
    );
  blk00000287_blk00000288_blk00000292 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000287_blk00000288_sig0000124d,
      Q => sig000002da
    );
  blk00000287_blk00000288_blk00000291 : SRLC32E
    generic map(
      INIT => X"00000000"
    )
    port map (
      CLK => clk,
      D => sig000002f4,
      CE => ce,
      Q => blk00000287_blk00000288_sig0000124d,
      Q31 => NLW_blk00000287_blk00000288_blk00000291_Q31_UNCONNECTED,
      A(4) => blk00000287_blk00000288_sig00001249,
      A(3) => blk00000287_blk00000288_sig00001249,
      A(2) => blk00000287_blk00000288_sig00001249,
      A(1) => blk00000287_blk00000288_sig00001248,
      A(0) => blk00000287_blk00000288_sig00001248
    );
  blk00000287_blk00000288_blk00000290 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000287_blk00000288_sig0000124c,
      Q => sig000002d9
    );
  blk00000287_blk00000288_blk0000028f : SRLC32E
    generic map(
      INIT => X"00000000"
    )
    port map (
      CLK => clk,
      D => sig000002f3,
      CE => ce,
      Q => blk00000287_blk00000288_sig0000124c,
      Q31 => NLW_blk00000287_blk00000288_blk0000028f_Q31_UNCONNECTED,
      A(4) => blk00000287_blk00000288_sig00001249,
      A(3) => blk00000287_blk00000288_sig00001249,
      A(2) => blk00000287_blk00000288_sig00001249,
      A(1) => blk00000287_blk00000288_sig00001248,
      A(0) => blk00000287_blk00000288_sig00001248
    );
  blk00000287_blk00000288_blk0000028e : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000287_blk00000288_sig0000124b,
      Q => sig000002d8
    );
  blk00000287_blk00000288_blk0000028d : SRLC32E
    generic map(
      INIT => X"00000000"
    )
    port map (
      CLK => clk,
      D => sig000002f2,
      CE => ce,
      Q => blk00000287_blk00000288_sig0000124b,
      Q31 => NLW_blk00000287_blk00000288_blk0000028d_Q31_UNCONNECTED,
      A(4) => blk00000287_blk00000288_sig00001249,
      A(3) => blk00000287_blk00000288_sig00001249,
      A(2) => blk00000287_blk00000288_sig00001249,
      A(1) => blk00000287_blk00000288_sig00001248,
      A(0) => blk00000287_blk00000288_sig00001248
    );
  blk00000287_blk00000288_blk0000028c : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000287_blk00000288_sig0000124a,
      Q => sig000002d7
    );
  blk00000287_blk00000288_blk0000028b : SRLC32E
    generic map(
      INIT => X"00000000"
    )
    port map (
      CLK => clk,
      D => sig000002f1,
      CE => ce,
      Q => blk00000287_blk00000288_sig0000124a,
      Q31 => NLW_blk00000287_blk00000288_blk0000028b_Q31_UNCONNECTED,
      A(4) => blk00000287_blk00000288_sig00001249,
      A(3) => blk00000287_blk00000288_sig00001249,
      A(2) => blk00000287_blk00000288_sig00001249,
      A(1) => blk00000287_blk00000288_sig00001248,
      A(0) => blk00000287_blk00000288_sig00001248
    );
  blk00000287_blk00000288_blk0000028a : VCC
    port map (
      P => blk00000287_blk00000288_sig00001249
    );
  blk00000287_blk00000288_blk00000289 : GND
    port map (
      G => blk00000287_blk00000288_sig00001248
    );
  blk000002bf_blk000002f7 : LUT3
    generic map(
      INIT => X"6A"
    )
    port map (
      I0 => sig000002f0,
      I1 => sig00000324,
      I2 => sig0000030c,
      O => blk000002bf_sig000012b8
    );
  blk000002bf_blk000002f6 : LUT3
    generic map(
      INIT => X"6A"
    )
    port map (
      I0 => sig000002ed,
      I1 => sig00000322,
      I2 => sig0000030c,
      O => blk000002bf_sig000012ae
    );
  blk000002bf_blk000002f5 : LUT3
    generic map(
      INIT => X"6A"
    )
    port map (
      I0 => sig000002ec,
      I1 => sig00000321,
      I2 => sig0000030c,
      O => blk000002bf_sig000012af
    );
  blk000002bf_blk000002f4 : LUT3
    generic map(
      INIT => X"6A"
    )
    port map (
      I0 => sig000002eb,
      I1 => sig00000320,
      I2 => sig0000030c,
      O => blk000002bf_sig000012b0
    );
  blk000002bf_blk000002f3 : LUT3
    generic map(
      INIT => X"6A"
    )
    port map (
      I0 => sig000002ea,
      I1 => sig0000031f,
      I2 => sig0000030c,
      O => blk000002bf_sig000012b1
    );
  blk000002bf_blk000002f2 : LUT3
    generic map(
      INIT => X"6A"
    )
    port map (
      I0 => sig000002e9,
      I1 => sig0000031e,
      I2 => sig0000030c,
      O => blk000002bf_sig000012b2
    );
  blk000002bf_blk000002f1 : LUT3
    generic map(
      INIT => X"6A"
    )
    port map (
      I0 => sig000002e8,
      I1 => sig0000031d,
      I2 => sig0000030c,
      O => blk000002bf_sig000012b3
    );
  blk000002bf_blk000002f0 : LUT3
    generic map(
      INIT => X"6A"
    )
    port map (
      I0 => sig000002e7,
      I1 => sig0000031c,
      I2 => sig0000030c,
      O => blk000002bf_sig000012b4
    );
  blk000002bf_blk000002ef : LUT3
    generic map(
      INIT => X"6A"
    )
    port map (
      I0 => sig000002e6,
      I1 => sig0000031b,
      I2 => sig0000030c,
      O => blk000002bf_sig000012b5
    );
  blk000002bf_blk000002ee : LUT3
    generic map(
      INIT => X"6A"
    )
    port map (
      I0 => sig000002e5,
      I1 => sig0000031a,
      I2 => sig0000030c,
      O => blk000002bf_sig000012b6
    );
  blk000002bf_blk000002ed : LUT3
    generic map(
      INIT => X"6A"
    )
    port map (
      I0 => sig000002f0,
      I1 => sig00000324,
      I2 => sig0000030c,
      O => blk000002bf_sig000012ab
    );
  blk000002bf_blk000002ec : LUT3
    generic map(
      INIT => X"6A"
    )
    port map (
      I0 => sig000002ef,
      I1 => sig00000324,
      I2 => sig0000030c,
      O => blk000002bf_sig000012ac
    );
  blk000002bf_blk000002eb : LUT3
    generic map(
      INIT => X"6A"
    )
    port map (
      I0 => sig000002ee,
      I1 => sig00000323,
      I2 => sig0000030c,
      O => blk000002bf_sig000012ad
    );
  blk000002bf_blk000002ea : LUT3
    generic map(
      INIT => X"6A"
    )
    port map (
      I0 => sig000002e4,
      I1 => sig00000319,
      I2 => sig0000030c,
      O => blk000002bf_sig000012b7
    );
  blk000002bf_blk000002e9 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk000002bf_sig000012a9,
      Q => sig0000026e
    );
  blk000002bf_blk000002e8 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk000002bf_sig0000129b,
      Q => sig0000026f
    );
  blk000002bf_blk000002e7 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk000002bf_sig0000129a,
      Q => sig00000270
    );
  blk000002bf_blk000002e6 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk000002bf_sig00001299,
      Q => sig00000271
    );
  blk000002bf_blk000002e5 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk000002bf_sig00001298,
      Q => sig00000272
    );
  blk000002bf_blk000002e4 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk000002bf_sig00001297,
      Q => sig00000273
    );
  blk000002bf_blk000002e3 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk000002bf_sig00001296,
      Q => sig00000274
    );
  blk000002bf_blk000002e2 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk000002bf_sig00001295,
      Q => sig00000275
    );
  blk000002bf_blk000002e1 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk000002bf_sig00001294,
      Q => sig00000276
    );
  blk000002bf_blk000002e0 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk000002bf_sig00001293,
      Q => sig00000277
    );
  blk000002bf_blk000002df : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk000002bf_sig00001292,
      Q => sig00000278
    );
  blk000002bf_blk000002de : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk000002bf_sig00001291,
      Q => sig00000279
    );
  blk000002bf_blk000002dd : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk000002bf_sig00001290,
      Q => sig0000027a
    );
  blk000002bf_blk000002dc : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk000002bf_sig0000129c,
      Q => sig000002b9
    );
  blk000002bf_blk000002db : MUXCY
    port map (
      CI => blk000002bf_sig0000128f,
      DI => sig000002e4,
      S => blk000002bf_sig000012b7,
      O => blk000002bf_sig000012aa
    );
  blk000002bf_blk000002da : XORCY
    port map (
      CI => blk000002bf_sig0000128f,
      LI => blk000002bf_sig000012b7,
      O => blk000002bf_sig000012a9
    );
  blk000002bf_blk000002d9 : MUXCY
    port map (
      CI => blk000002bf_sig000012aa,
      DI => sig000002e5,
      S => blk000002bf_sig000012b6,
      O => blk000002bf_sig000012a8
    );
  blk000002bf_blk000002d8 : MUXCY
    port map (
      CI => blk000002bf_sig000012a8,
      DI => sig000002e6,
      S => blk000002bf_sig000012b5,
      O => blk000002bf_sig000012a7
    );
  blk000002bf_blk000002d7 : MUXCY
    port map (
      CI => blk000002bf_sig000012a7,
      DI => sig000002e7,
      S => blk000002bf_sig000012b4,
      O => blk000002bf_sig000012a6
    );
  blk000002bf_blk000002d6 : MUXCY
    port map (
      CI => blk000002bf_sig000012a6,
      DI => sig000002e8,
      S => blk000002bf_sig000012b3,
      O => blk000002bf_sig000012a5
    );
  blk000002bf_blk000002d5 : MUXCY
    port map (
      CI => blk000002bf_sig000012a5,
      DI => sig000002e9,
      S => blk000002bf_sig000012b2,
      O => blk000002bf_sig000012a4
    );
  blk000002bf_blk000002d4 : MUXCY
    port map (
      CI => blk000002bf_sig000012a4,
      DI => sig000002ea,
      S => blk000002bf_sig000012b1,
      O => blk000002bf_sig000012a3
    );
  blk000002bf_blk000002d3 : MUXCY
    port map (
      CI => blk000002bf_sig000012a3,
      DI => sig000002eb,
      S => blk000002bf_sig000012b0,
      O => blk000002bf_sig000012a2
    );
  blk000002bf_blk000002d2 : MUXCY
    port map (
      CI => blk000002bf_sig000012a2,
      DI => sig000002ec,
      S => blk000002bf_sig000012af,
      O => blk000002bf_sig000012a1
    );
  blk000002bf_blk000002d1 : MUXCY
    port map (
      CI => blk000002bf_sig000012a1,
      DI => sig000002ed,
      S => blk000002bf_sig000012ae,
      O => blk000002bf_sig000012a0
    );
  blk000002bf_blk000002d0 : MUXCY
    port map (
      CI => blk000002bf_sig000012a0,
      DI => sig000002ee,
      S => blk000002bf_sig000012ad,
      O => blk000002bf_sig0000129f
    );
  blk000002bf_blk000002cf : MUXCY
    port map (
      CI => blk000002bf_sig0000129f,
      DI => sig000002ef,
      S => blk000002bf_sig000012ac,
      O => blk000002bf_sig0000129e
    );
  blk000002bf_blk000002ce : MUXCY
    port map (
      CI => blk000002bf_sig0000129e,
      DI => sig000002f0,
      S => blk000002bf_sig000012b8,
      O => blk000002bf_sig0000129d
    );
  blk000002bf_blk000002cd : XORCY
    port map (
      CI => blk000002bf_sig0000129d,
      LI => blk000002bf_sig000012ab,
      O => blk000002bf_sig0000129c
    );
  blk000002bf_blk000002cc : XORCY
    port map (
      CI => blk000002bf_sig000012aa,
      LI => blk000002bf_sig000012b6,
      O => blk000002bf_sig0000129b
    );
  blk000002bf_blk000002cb : XORCY
    port map (
      CI => blk000002bf_sig000012a8,
      LI => blk000002bf_sig000012b5,
      O => blk000002bf_sig0000129a
    );
  blk000002bf_blk000002ca : XORCY
    port map (
      CI => blk000002bf_sig000012a7,
      LI => blk000002bf_sig000012b4,
      O => blk000002bf_sig00001299
    );
  blk000002bf_blk000002c9 : XORCY
    port map (
      CI => blk000002bf_sig000012a6,
      LI => blk000002bf_sig000012b3,
      O => blk000002bf_sig00001298
    );
  blk000002bf_blk000002c8 : XORCY
    port map (
      CI => blk000002bf_sig000012a5,
      LI => blk000002bf_sig000012b2,
      O => blk000002bf_sig00001297
    );
  blk000002bf_blk000002c7 : XORCY
    port map (
      CI => blk000002bf_sig000012a4,
      LI => blk000002bf_sig000012b1,
      O => blk000002bf_sig00001296
    );
  blk000002bf_blk000002c6 : XORCY
    port map (
      CI => blk000002bf_sig000012a3,
      LI => blk000002bf_sig000012b0,
      O => blk000002bf_sig00001295
    );
  blk000002bf_blk000002c5 : XORCY
    port map (
      CI => blk000002bf_sig000012a2,
      LI => blk000002bf_sig000012af,
      O => blk000002bf_sig00001294
    );
  blk000002bf_blk000002c4 : XORCY
    port map (
      CI => blk000002bf_sig000012a1,
      LI => blk000002bf_sig000012ae,
      O => blk000002bf_sig00001293
    );
  blk000002bf_blk000002c3 : XORCY
    port map (
      CI => blk000002bf_sig000012a0,
      LI => blk000002bf_sig000012ad,
      O => blk000002bf_sig00001292
    );
  blk000002bf_blk000002c2 : XORCY
    port map (
      CI => blk000002bf_sig0000129f,
      LI => blk000002bf_sig000012ac,
      O => blk000002bf_sig00001291
    );
  blk000002bf_blk000002c1 : XORCY
    port map (
      CI => blk000002bf_sig0000129e,
      LI => blk000002bf_sig000012b8,
      O => blk000002bf_sig00001290
    );
  blk000002bf_blk000002c0 : GND
    port map (
      G => blk000002bf_sig0000128f
    );
  blk000002f8_blk00000330 : LUT3
    generic map(
      INIT => X"6A"
    )
    port map (
      I0 => sig000002e3,
      I1 => sig00000318,
      I2 => sig0000030c,
      O => blk000002f8_sig0000130d
    );
  blk000002f8_blk0000032f : LUT3
    generic map(
      INIT => X"6A"
    )
    port map (
      I0 => sig000002e0,
      I1 => sig00000316,
      I2 => sig0000030c,
      O => blk000002f8_sig00001303
    );
  blk000002f8_blk0000032e : LUT3
    generic map(
      INIT => X"6A"
    )
    port map (
      I0 => sig000002df,
      I1 => sig00000315,
      I2 => sig0000030c,
      O => blk000002f8_sig00001304
    );
  blk000002f8_blk0000032d : LUT3
    generic map(
      INIT => X"6A"
    )
    port map (
      I0 => sig000002de,
      I1 => sig00000314,
      I2 => sig0000030c,
      O => blk000002f8_sig00001305
    );
  blk000002f8_blk0000032c : LUT3
    generic map(
      INIT => X"6A"
    )
    port map (
      I0 => sig000002dd,
      I1 => sig00000313,
      I2 => sig0000030c,
      O => blk000002f8_sig00001306
    );
  blk000002f8_blk0000032b : LUT3
    generic map(
      INIT => X"6A"
    )
    port map (
      I0 => sig000002dc,
      I1 => sig00000312,
      I2 => sig0000030c,
      O => blk000002f8_sig00001307
    );
  blk000002f8_blk0000032a : LUT3
    generic map(
      INIT => X"6A"
    )
    port map (
      I0 => sig000002db,
      I1 => sig00000311,
      I2 => sig0000030c,
      O => blk000002f8_sig00001308
    );
  blk000002f8_blk00000329 : LUT3
    generic map(
      INIT => X"6A"
    )
    port map (
      I0 => sig000002da,
      I1 => sig00000310,
      I2 => sig0000030c,
      O => blk000002f8_sig00001309
    );
  blk000002f8_blk00000328 : LUT3
    generic map(
      INIT => X"6A"
    )
    port map (
      I0 => sig000002d9,
      I1 => sig0000030f,
      I2 => sig0000030c,
      O => blk000002f8_sig0000130a
    );
  blk000002f8_blk00000327 : LUT3
    generic map(
      INIT => X"6A"
    )
    port map (
      I0 => sig000002d8,
      I1 => sig0000030e,
      I2 => sig0000030c,
      O => blk000002f8_sig0000130b
    );
  blk000002f8_blk00000326 : LUT3
    generic map(
      INIT => X"6A"
    )
    port map (
      I0 => sig000002e3,
      I1 => sig00000318,
      I2 => sig0000030c,
      O => blk000002f8_sig00001300
    );
  blk000002f8_blk00000325 : LUT3
    generic map(
      INIT => X"6A"
    )
    port map (
      I0 => sig000002e2,
      I1 => sig00000318,
      I2 => sig0000030c,
      O => blk000002f8_sig00001301
    );
  blk000002f8_blk00000324 : LUT3
    generic map(
      INIT => X"6A"
    )
    port map (
      I0 => sig000002e1,
      I1 => sig00000317,
      I2 => sig0000030c,
      O => blk000002f8_sig00001302
    );
  blk000002f8_blk00000323 : LUT3
    generic map(
      INIT => X"6A"
    )
    port map (
      I0 => sig000002d7,
      I1 => sig0000030d,
      I2 => sig0000030c,
      O => blk000002f8_sig0000130c
    );
  blk000002f8_blk00000322 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk000002f8_sig000012fe,
      Q => sig00000261
    );
  blk000002f8_blk00000321 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk000002f8_sig000012f0,
      Q => sig00000262
    );
  blk000002f8_blk00000320 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk000002f8_sig000012ef,
      Q => sig00000263
    );
  blk000002f8_blk0000031f : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk000002f8_sig000012ee,
      Q => sig00000264
    );
  blk000002f8_blk0000031e : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk000002f8_sig000012ed,
      Q => sig00000265
    );
  blk000002f8_blk0000031d : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk000002f8_sig000012ec,
      Q => sig00000266
    );
  blk000002f8_blk0000031c : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk000002f8_sig000012eb,
      Q => sig00000267
    );
  blk000002f8_blk0000031b : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk000002f8_sig000012ea,
      Q => sig00000268
    );
  blk000002f8_blk0000031a : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk000002f8_sig000012e9,
      Q => sig00000269
    );
  blk000002f8_blk00000319 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk000002f8_sig000012e8,
      Q => sig0000026a
    );
  blk000002f8_blk00000318 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk000002f8_sig000012e7,
      Q => sig0000026b
    );
  blk000002f8_blk00000317 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk000002f8_sig000012e6,
      Q => sig0000026c
    );
  blk000002f8_blk00000316 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk000002f8_sig000012e5,
      Q => sig0000026d
    );
  blk000002f8_blk00000315 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk000002f8_sig000012f1,
      Q => sig000002bb
    );
  blk000002f8_blk00000314 : MUXCY
    port map (
      CI => blk000002f8_sig000012e4,
      DI => sig000002d7,
      S => blk000002f8_sig0000130c,
      O => blk000002f8_sig000012ff
    );
  blk000002f8_blk00000313 : XORCY
    port map (
      CI => blk000002f8_sig000012e4,
      LI => blk000002f8_sig0000130c,
      O => blk000002f8_sig000012fe
    );
  blk000002f8_blk00000312 : MUXCY
    port map (
      CI => blk000002f8_sig000012ff,
      DI => sig000002d8,
      S => blk000002f8_sig0000130b,
      O => blk000002f8_sig000012fd
    );
  blk000002f8_blk00000311 : MUXCY
    port map (
      CI => blk000002f8_sig000012fd,
      DI => sig000002d9,
      S => blk000002f8_sig0000130a,
      O => blk000002f8_sig000012fc
    );
  blk000002f8_blk00000310 : MUXCY
    port map (
      CI => blk000002f8_sig000012fc,
      DI => sig000002da,
      S => blk000002f8_sig00001309,
      O => blk000002f8_sig000012fb
    );
  blk000002f8_blk0000030f : MUXCY
    port map (
      CI => blk000002f8_sig000012fb,
      DI => sig000002db,
      S => blk000002f8_sig00001308,
      O => blk000002f8_sig000012fa
    );
  blk000002f8_blk0000030e : MUXCY
    port map (
      CI => blk000002f8_sig000012fa,
      DI => sig000002dc,
      S => blk000002f8_sig00001307,
      O => blk000002f8_sig000012f9
    );
  blk000002f8_blk0000030d : MUXCY
    port map (
      CI => blk000002f8_sig000012f9,
      DI => sig000002dd,
      S => blk000002f8_sig00001306,
      O => blk000002f8_sig000012f8
    );
  blk000002f8_blk0000030c : MUXCY
    port map (
      CI => blk000002f8_sig000012f8,
      DI => sig000002de,
      S => blk000002f8_sig00001305,
      O => blk000002f8_sig000012f7
    );
  blk000002f8_blk0000030b : MUXCY
    port map (
      CI => blk000002f8_sig000012f7,
      DI => sig000002df,
      S => blk000002f8_sig00001304,
      O => blk000002f8_sig000012f6
    );
  blk000002f8_blk0000030a : MUXCY
    port map (
      CI => blk000002f8_sig000012f6,
      DI => sig000002e0,
      S => blk000002f8_sig00001303,
      O => blk000002f8_sig000012f5
    );
  blk000002f8_blk00000309 : MUXCY
    port map (
      CI => blk000002f8_sig000012f5,
      DI => sig000002e1,
      S => blk000002f8_sig00001302,
      O => blk000002f8_sig000012f4
    );
  blk000002f8_blk00000308 : MUXCY
    port map (
      CI => blk000002f8_sig000012f4,
      DI => sig000002e2,
      S => blk000002f8_sig00001301,
      O => blk000002f8_sig000012f3
    );
  blk000002f8_blk00000307 : MUXCY
    port map (
      CI => blk000002f8_sig000012f3,
      DI => sig000002e3,
      S => blk000002f8_sig0000130d,
      O => blk000002f8_sig000012f2
    );
  blk000002f8_blk00000306 : XORCY
    port map (
      CI => blk000002f8_sig000012f2,
      LI => blk000002f8_sig00001300,
      O => blk000002f8_sig000012f1
    );
  blk000002f8_blk00000305 : XORCY
    port map (
      CI => blk000002f8_sig000012ff,
      LI => blk000002f8_sig0000130b,
      O => blk000002f8_sig000012f0
    );
  blk000002f8_blk00000304 : XORCY
    port map (
      CI => blk000002f8_sig000012fd,
      LI => blk000002f8_sig0000130a,
      O => blk000002f8_sig000012ef
    );
  blk000002f8_blk00000303 : XORCY
    port map (
      CI => blk000002f8_sig000012fc,
      LI => blk000002f8_sig00001309,
      O => blk000002f8_sig000012ee
    );
  blk000002f8_blk00000302 : XORCY
    port map (
      CI => blk000002f8_sig000012fb,
      LI => blk000002f8_sig00001308,
      O => blk000002f8_sig000012ed
    );
  blk000002f8_blk00000301 : XORCY
    port map (
      CI => blk000002f8_sig000012fa,
      LI => blk000002f8_sig00001307,
      O => blk000002f8_sig000012ec
    );
  blk000002f8_blk00000300 : XORCY
    port map (
      CI => blk000002f8_sig000012f9,
      LI => blk000002f8_sig00001306,
      O => blk000002f8_sig000012eb
    );
  blk000002f8_blk000002ff : XORCY
    port map (
      CI => blk000002f8_sig000012f8,
      LI => blk000002f8_sig00001305,
      O => blk000002f8_sig000012ea
    );
  blk000002f8_blk000002fe : XORCY
    port map (
      CI => blk000002f8_sig000012f7,
      LI => blk000002f8_sig00001304,
      O => blk000002f8_sig000012e9
    );
  blk000002f8_blk000002fd : XORCY
    port map (
      CI => blk000002f8_sig000012f6,
      LI => blk000002f8_sig00001303,
      O => blk000002f8_sig000012e8
    );
  blk000002f8_blk000002fc : XORCY
    port map (
      CI => blk000002f8_sig000012f5,
      LI => blk000002f8_sig00001302,
      O => blk000002f8_sig000012e7
    );
  blk000002f8_blk000002fb : XORCY
    port map (
      CI => blk000002f8_sig000012f4,
      LI => blk000002f8_sig00001301,
      O => blk000002f8_sig000012e6
    );
  blk000002f8_blk000002fa : XORCY
    port map (
      CI => blk000002f8_sig000012f3,
      LI => blk000002f8_sig0000130d,
      O => blk000002f8_sig000012e5
    );
  blk000002f8_blk000002f9 : GND
    port map (
      G => blk000002f8_sig000012e4
    );
  blk00000331_blk00000375 : LUT3
    generic map(
      INIT => X"9A"
    )
    port map (
      I0 => sig00000324,
      I1 => sig000002f0,
      I2 => sig0000030c,
      O => blk00000331_sig0000136e
    );
  blk00000331_blk00000374 : LUT2
    generic map(
      INIT => X"8"
    )
    port map (
      I0 => sig000002e4,
      I1 => sig0000030c,
      O => blk00000331_sig0000135c
    );
  blk00000331_blk00000373 : LUT2
    generic map(
      INIT => X"8"
    )
    port map (
      I0 => sig000002e5,
      I1 => sig0000030c,
      O => blk00000331_sig0000135b
    );
  blk00000331_blk00000372 : LUT2
    generic map(
      INIT => X"8"
    )
    port map (
      I0 => sig000002e6,
      I1 => sig0000030c,
      O => blk00000331_sig0000135a
    );
  blk00000331_blk00000371 : LUT2
    generic map(
      INIT => X"8"
    )
    port map (
      I0 => sig000002e7,
      I1 => sig0000030c,
      O => blk00000331_sig00001359
    );
  blk00000331_blk00000370 : LUT2
    generic map(
      INIT => X"8"
    )
    port map (
      I0 => sig000002e8,
      I1 => sig0000030c,
      O => blk00000331_sig00001358
    );
  blk00000331_blk0000036f : LUT2
    generic map(
      INIT => X"8"
    )
    port map (
      I0 => sig000002e9,
      I1 => sig0000030c,
      O => blk00000331_sig00001357
    );
  blk00000331_blk0000036e : LUT2
    generic map(
      INIT => X"8"
    )
    port map (
      I0 => sig000002ea,
      I1 => sig0000030c,
      O => blk00000331_sig00001356
    );
  blk00000331_blk0000036d : LUT2
    generic map(
      INIT => X"8"
    )
    port map (
      I0 => sig000002eb,
      I1 => sig0000030c,
      O => blk00000331_sig00001355
    );
  blk00000331_blk0000036c : LUT2
    generic map(
      INIT => X"8"
    )
    port map (
      I0 => sig000002ec,
      I1 => sig0000030c,
      O => blk00000331_sig00001354
    );
  blk00000331_blk0000036b : LUT2
    generic map(
      INIT => X"8"
    )
    port map (
      I0 => sig000002ed,
      I1 => sig0000030c,
      O => blk00000331_sig00001353
    );
  blk00000331_blk0000036a : LUT2
    generic map(
      INIT => X"8"
    )
    port map (
      I0 => sig000002ee,
      I1 => sig0000030c,
      O => blk00000331_sig00001352
    );
  blk00000331_blk00000369 : LUT2
    generic map(
      INIT => X"8"
    )
    port map (
      I0 => sig000002ef,
      I1 => sig0000030c,
      O => blk00000331_sig00001351
    );
  blk00000331_blk00000368 : LUT2
    generic map(
      INIT => X"8"
    )
    port map (
      I0 => sig000002f0,
      I1 => sig0000030c,
      O => blk00000331_sig00001350
    );
  blk00000331_blk00000367 : LUT3
    generic map(
      INIT => X"9A"
    )
    port map (
      I0 => sig00000322,
      I1 => sig000002ed,
      I2 => sig0000030c,
      O => blk00000331_sig00001364
    );
  blk00000331_blk00000366 : LUT3
    generic map(
      INIT => X"9A"
    )
    port map (
      I0 => sig00000321,
      I1 => sig000002ec,
      I2 => sig0000030c,
      O => blk00000331_sig00001365
    );
  blk00000331_blk00000365 : LUT3
    generic map(
      INIT => X"9A"
    )
    port map (
      I0 => sig00000320,
      I1 => sig000002eb,
      I2 => sig0000030c,
      O => blk00000331_sig00001366
    );
  blk00000331_blk00000364 : LUT3
    generic map(
      INIT => X"9A"
    )
    port map (
      I0 => sig0000031f,
      I1 => sig000002ea,
      I2 => sig0000030c,
      O => blk00000331_sig00001367
    );
  blk00000331_blk00000363 : LUT3
    generic map(
      INIT => X"9A"
    )
    port map (
      I0 => sig0000031e,
      I1 => sig000002e9,
      I2 => sig0000030c,
      O => blk00000331_sig00001368
    );
  blk00000331_blk00000362 : LUT3
    generic map(
      INIT => X"9A"
    )
    port map (
      I0 => sig0000031d,
      I1 => sig000002e8,
      I2 => sig0000030c,
      O => blk00000331_sig00001369
    );
  blk00000331_blk00000361 : LUT3
    generic map(
      INIT => X"9A"
    )
    port map (
      I0 => sig0000031c,
      I1 => sig000002e7,
      I2 => sig0000030c,
      O => blk00000331_sig0000136a
    );
  blk00000331_blk00000360 : LUT3
    generic map(
      INIT => X"9A"
    )
    port map (
      I0 => sig0000031b,
      I1 => sig000002e6,
      I2 => sig0000030c,
      O => blk00000331_sig0000136b
    );
  blk00000331_blk0000035f : LUT3
    generic map(
      INIT => X"9A"
    )
    port map (
      I0 => sig0000031a,
      I1 => sig000002e5,
      I2 => sig0000030c,
      O => blk00000331_sig0000136c
    );
  blk00000331_blk0000035e : LUT3
    generic map(
      INIT => X"9A"
    )
    port map (
      I0 => sig00000324,
      I1 => sig000002f0,
      I2 => sig0000030c,
      O => blk00000331_sig00001361
    );
  blk00000331_blk0000035d : LUT3
    generic map(
      INIT => X"9A"
    )
    port map (
      I0 => sig00000324,
      I1 => sig000002ef,
      I2 => sig0000030c,
      O => blk00000331_sig00001362
    );
  blk00000331_blk0000035c : LUT3
    generic map(
      INIT => X"9A"
    )
    port map (
      I0 => sig00000323,
      I1 => sig000002ee,
      I2 => sig0000030c,
      O => blk00000331_sig00001363
    );
  blk00000331_blk0000035b : LUT3
    generic map(
      INIT => X"9A"
    )
    port map (
      I0 => sig00000319,
      I1 => sig000002e4,
      I2 => sig0000030c,
      O => blk00000331_sig0000136d
    );
  blk00000331_blk0000035a : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000331_sig0000135f,
      Q => sig000002ca
    );
  blk00000331_blk00000359 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000331_sig0000135d,
      Q => sig000002cb
    );
  blk00000331_blk00000358 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000331_sig0000134d,
      Q => sig000002cc
    );
  blk00000331_blk00000357 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000331_sig0000134b,
      Q => sig000002cd
    );
  blk00000331_blk00000356 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000331_sig00001349,
      Q => sig000002ce
    );
  blk00000331_blk00000355 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000331_sig00001347,
      Q => sig000002cf
    );
  blk00000331_blk00000354 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000331_sig00001345,
      Q => sig000002d0
    );
  blk00000331_blk00000353 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000331_sig00001343,
      Q => sig000002d1
    );
  blk00000331_blk00000352 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000331_sig00001341,
      Q => sig000002d2
    );
  blk00000331_blk00000351 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000331_sig0000133f,
      Q => sig000002d3
    );
  blk00000331_blk00000350 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000331_sig0000133d,
      Q => sig000002d4
    );
  blk00000331_blk0000034f : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000331_sig0000133b,
      Q => sig000002d5
    );
  blk00000331_blk0000034e : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000331_sig00001339,
      Q => sig000002d6
    );
  blk00000331_blk0000034d : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000331_sig0000134f,
      Q => sig000002ba
    );
  blk00000331_blk0000034c : MUXCY
    port map (
      CI => sig0000030c,
      DI => blk00000331_sig0000135c,
      S => blk00000331_sig0000136d,
      O => blk00000331_sig00001360
    );
  blk00000331_blk0000034b : XORCY
    port map (
      CI => sig0000030c,
      LI => blk00000331_sig0000136d,
      O => blk00000331_sig0000135f
    );
  blk00000331_blk0000034a : MUXCY
    port map (
      CI => blk00000331_sig00001360,
      DI => blk00000331_sig0000135b,
      S => blk00000331_sig0000136c,
      O => blk00000331_sig0000135e
    );
  blk00000331_blk00000349 : XORCY
    port map (
      CI => blk00000331_sig00001360,
      LI => blk00000331_sig0000136c,
      O => blk00000331_sig0000135d
    );
  blk00000331_blk00000348 : XORCY
    port map (
      CI => blk00000331_sig0000133a,
      LI => blk00000331_sig00001361,
      O => blk00000331_sig0000134f
    );
  blk00000331_blk00000347 : MUXCY
    port map (
      CI => blk00000331_sig0000135e,
      DI => blk00000331_sig0000135a,
      S => blk00000331_sig0000136b,
      O => blk00000331_sig0000134e
    );
  blk00000331_blk00000346 : XORCY
    port map (
      CI => blk00000331_sig0000135e,
      LI => blk00000331_sig0000136b,
      O => blk00000331_sig0000134d
    );
  blk00000331_blk00000345 : MUXCY
    port map (
      CI => blk00000331_sig0000134e,
      DI => blk00000331_sig00001359,
      S => blk00000331_sig0000136a,
      O => blk00000331_sig0000134c
    );
  blk00000331_blk00000344 : XORCY
    port map (
      CI => blk00000331_sig0000134e,
      LI => blk00000331_sig0000136a,
      O => blk00000331_sig0000134b
    );
  blk00000331_blk00000343 : MUXCY
    port map (
      CI => blk00000331_sig0000134c,
      DI => blk00000331_sig00001358,
      S => blk00000331_sig00001369,
      O => blk00000331_sig0000134a
    );
  blk00000331_blk00000342 : XORCY
    port map (
      CI => blk00000331_sig0000134c,
      LI => blk00000331_sig00001369,
      O => blk00000331_sig00001349
    );
  blk00000331_blk00000341 : MUXCY
    port map (
      CI => blk00000331_sig0000134a,
      DI => blk00000331_sig00001357,
      S => blk00000331_sig00001368,
      O => blk00000331_sig00001348
    );
  blk00000331_blk00000340 : XORCY
    port map (
      CI => blk00000331_sig0000134a,
      LI => blk00000331_sig00001368,
      O => blk00000331_sig00001347
    );
  blk00000331_blk0000033f : MUXCY
    port map (
      CI => blk00000331_sig00001348,
      DI => blk00000331_sig00001356,
      S => blk00000331_sig00001367,
      O => blk00000331_sig00001346
    );
  blk00000331_blk0000033e : XORCY
    port map (
      CI => blk00000331_sig00001348,
      LI => blk00000331_sig00001367,
      O => blk00000331_sig00001345
    );
  blk00000331_blk0000033d : MUXCY
    port map (
      CI => blk00000331_sig00001346,
      DI => blk00000331_sig00001355,
      S => blk00000331_sig00001366,
      O => blk00000331_sig00001344
    );
  blk00000331_blk0000033c : XORCY
    port map (
      CI => blk00000331_sig00001346,
      LI => blk00000331_sig00001366,
      O => blk00000331_sig00001343
    );
  blk00000331_blk0000033b : MUXCY
    port map (
      CI => blk00000331_sig00001344,
      DI => blk00000331_sig00001354,
      S => blk00000331_sig00001365,
      O => blk00000331_sig00001342
    );
  blk00000331_blk0000033a : XORCY
    port map (
      CI => blk00000331_sig00001344,
      LI => blk00000331_sig00001365,
      O => blk00000331_sig00001341
    );
  blk00000331_blk00000339 : MUXCY
    port map (
      CI => blk00000331_sig00001342,
      DI => blk00000331_sig00001353,
      S => blk00000331_sig00001364,
      O => blk00000331_sig00001340
    );
  blk00000331_blk00000338 : XORCY
    port map (
      CI => blk00000331_sig00001342,
      LI => blk00000331_sig00001364,
      O => blk00000331_sig0000133f
    );
  blk00000331_blk00000337 : MUXCY
    port map (
      CI => blk00000331_sig00001340,
      DI => blk00000331_sig00001352,
      S => blk00000331_sig00001363,
      O => blk00000331_sig0000133e
    );
  blk00000331_blk00000336 : XORCY
    port map (
      CI => blk00000331_sig00001340,
      LI => blk00000331_sig00001363,
      O => blk00000331_sig0000133d
    );
  blk00000331_blk00000335 : MUXCY
    port map (
      CI => blk00000331_sig0000133e,
      DI => blk00000331_sig00001351,
      S => blk00000331_sig00001362,
      O => blk00000331_sig0000133c
    );
  blk00000331_blk00000334 : XORCY
    port map (
      CI => blk00000331_sig0000133e,
      LI => blk00000331_sig00001362,
      O => blk00000331_sig0000133b
    );
  blk00000331_blk00000333 : MUXCY
    port map (
      CI => blk00000331_sig0000133c,
      DI => blk00000331_sig00001350,
      S => blk00000331_sig0000136e,
      O => blk00000331_sig0000133a
    );
  blk00000331_blk00000332 : XORCY
    port map (
      CI => blk00000331_sig0000133c,
      LI => blk00000331_sig0000136e,
      O => blk00000331_sig00001339
    );
  blk00000376_blk000003ba : LUT3
    generic map(
      INIT => X"9A"
    )
    port map (
      I0 => sig00000318,
      I1 => sig000002e3,
      I2 => sig0000030c,
      O => blk00000376_sig000013cf
    );
  blk00000376_blk000003b9 : LUT2
    generic map(
      INIT => X"8"
    )
    port map (
      I0 => sig000002d7,
      I1 => sig0000030c,
      O => blk00000376_sig000013bd
    );
  blk00000376_blk000003b8 : LUT2
    generic map(
      INIT => X"8"
    )
    port map (
      I0 => sig000002d8,
      I1 => sig0000030c,
      O => blk00000376_sig000013bc
    );
  blk00000376_blk000003b7 : LUT2
    generic map(
      INIT => X"8"
    )
    port map (
      I0 => sig000002d9,
      I1 => sig0000030c,
      O => blk00000376_sig000013bb
    );
  blk00000376_blk000003b6 : LUT2
    generic map(
      INIT => X"8"
    )
    port map (
      I0 => sig000002da,
      I1 => sig0000030c,
      O => blk00000376_sig000013ba
    );
  blk00000376_blk000003b5 : LUT2
    generic map(
      INIT => X"8"
    )
    port map (
      I0 => sig000002db,
      I1 => sig0000030c,
      O => blk00000376_sig000013b9
    );
  blk00000376_blk000003b4 : LUT2
    generic map(
      INIT => X"8"
    )
    port map (
      I0 => sig000002dc,
      I1 => sig0000030c,
      O => blk00000376_sig000013b8
    );
  blk00000376_blk000003b3 : LUT2
    generic map(
      INIT => X"8"
    )
    port map (
      I0 => sig000002dd,
      I1 => sig0000030c,
      O => blk00000376_sig000013b7
    );
  blk00000376_blk000003b2 : LUT2
    generic map(
      INIT => X"8"
    )
    port map (
      I0 => sig000002de,
      I1 => sig0000030c,
      O => blk00000376_sig000013b6
    );
  blk00000376_blk000003b1 : LUT2
    generic map(
      INIT => X"8"
    )
    port map (
      I0 => sig000002df,
      I1 => sig0000030c,
      O => blk00000376_sig000013b5
    );
  blk00000376_blk000003b0 : LUT2
    generic map(
      INIT => X"8"
    )
    port map (
      I0 => sig000002e0,
      I1 => sig0000030c,
      O => blk00000376_sig000013b4
    );
  blk00000376_blk000003af : LUT2
    generic map(
      INIT => X"8"
    )
    port map (
      I0 => sig000002e1,
      I1 => sig0000030c,
      O => blk00000376_sig000013b3
    );
  blk00000376_blk000003ae : LUT2
    generic map(
      INIT => X"8"
    )
    port map (
      I0 => sig000002e2,
      I1 => sig0000030c,
      O => blk00000376_sig000013b2
    );
  blk00000376_blk000003ad : LUT2
    generic map(
      INIT => X"8"
    )
    port map (
      I0 => sig000002e3,
      I1 => sig0000030c,
      O => blk00000376_sig000013b1
    );
  blk00000376_blk000003ac : LUT3
    generic map(
      INIT => X"9A"
    )
    port map (
      I0 => sig00000316,
      I1 => sig000002e0,
      I2 => sig0000030c,
      O => blk00000376_sig000013c5
    );
  blk00000376_blk000003ab : LUT3
    generic map(
      INIT => X"9A"
    )
    port map (
      I0 => sig00000315,
      I1 => sig000002df,
      I2 => sig0000030c,
      O => blk00000376_sig000013c6
    );
  blk00000376_blk000003aa : LUT3
    generic map(
      INIT => X"9A"
    )
    port map (
      I0 => sig00000314,
      I1 => sig000002de,
      I2 => sig0000030c,
      O => blk00000376_sig000013c7
    );
  blk00000376_blk000003a9 : LUT3
    generic map(
      INIT => X"9A"
    )
    port map (
      I0 => sig00000313,
      I1 => sig000002dd,
      I2 => sig0000030c,
      O => blk00000376_sig000013c8
    );
  blk00000376_blk000003a8 : LUT3
    generic map(
      INIT => X"9A"
    )
    port map (
      I0 => sig00000312,
      I1 => sig000002dc,
      I2 => sig0000030c,
      O => blk00000376_sig000013c9
    );
  blk00000376_blk000003a7 : LUT3
    generic map(
      INIT => X"9A"
    )
    port map (
      I0 => sig00000311,
      I1 => sig000002db,
      I2 => sig0000030c,
      O => blk00000376_sig000013ca
    );
  blk00000376_blk000003a6 : LUT3
    generic map(
      INIT => X"9A"
    )
    port map (
      I0 => sig00000310,
      I1 => sig000002da,
      I2 => sig0000030c,
      O => blk00000376_sig000013cb
    );
  blk00000376_blk000003a5 : LUT3
    generic map(
      INIT => X"9A"
    )
    port map (
      I0 => sig0000030f,
      I1 => sig000002d9,
      I2 => sig0000030c,
      O => blk00000376_sig000013cc
    );
  blk00000376_blk000003a4 : LUT3
    generic map(
      INIT => X"9A"
    )
    port map (
      I0 => sig0000030e,
      I1 => sig000002d8,
      I2 => sig0000030c,
      O => blk00000376_sig000013cd
    );
  blk00000376_blk000003a3 : LUT3
    generic map(
      INIT => X"9A"
    )
    port map (
      I0 => sig00000318,
      I1 => sig000002e3,
      I2 => sig0000030c,
      O => blk00000376_sig000013c2
    );
  blk00000376_blk000003a2 : LUT3
    generic map(
      INIT => X"9A"
    )
    port map (
      I0 => sig00000318,
      I1 => sig000002e2,
      I2 => sig0000030c,
      O => blk00000376_sig000013c3
    );
  blk00000376_blk000003a1 : LUT3
    generic map(
      INIT => X"9A"
    )
    port map (
      I0 => sig00000317,
      I1 => sig000002e1,
      I2 => sig0000030c,
      O => blk00000376_sig000013c4
    );
  blk00000376_blk000003a0 : LUT3
    generic map(
      INIT => X"9A"
    )
    port map (
      I0 => sig0000030d,
      I1 => sig000002d7,
      I2 => sig0000030c,
      O => blk00000376_sig000013ce
    );
  blk00000376_blk0000039f : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000376_sig000013c0,
      Q => sig000002bd
    );
  blk00000376_blk0000039e : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000376_sig000013be,
      Q => sig000002be
    );
  blk00000376_blk0000039d : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000376_sig000013ae,
      Q => sig000002bf
    );
  blk00000376_blk0000039c : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000376_sig000013ac,
      Q => sig000002c0
    );
  blk00000376_blk0000039b : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000376_sig000013aa,
      Q => sig000002c1
    );
  blk00000376_blk0000039a : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000376_sig000013a8,
      Q => sig000002c2
    );
  blk00000376_blk00000399 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000376_sig000013a6,
      Q => sig000002c3
    );
  blk00000376_blk00000398 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000376_sig000013a4,
      Q => sig000002c4
    );
  blk00000376_blk00000397 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000376_sig000013a2,
      Q => sig000002c5
    );
  blk00000376_blk00000396 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000376_sig000013a0,
      Q => sig000002c6
    );
  blk00000376_blk00000395 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000376_sig0000139e,
      Q => sig000002c7
    );
  blk00000376_blk00000394 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000376_sig0000139c,
      Q => sig000002c8
    );
  blk00000376_blk00000393 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000376_sig0000139a,
      Q => sig000002c9
    );
  blk00000376_blk00000392 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000376_sig000013b0,
      Q => sig000002bc
    );
  blk00000376_blk00000391 : MUXCY
    port map (
      CI => sig0000030c,
      DI => blk00000376_sig000013bd,
      S => blk00000376_sig000013ce,
      O => blk00000376_sig000013c1
    );
  blk00000376_blk00000390 : XORCY
    port map (
      CI => sig0000030c,
      LI => blk00000376_sig000013ce,
      O => blk00000376_sig000013c0
    );
  blk00000376_blk0000038f : MUXCY
    port map (
      CI => blk00000376_sig000013c1,
      DI => blk00000376_sig000013bc,
      S => blk00000376_sig000013cd,
      O => blk00000376_sig000013bf
    );
  blk00000376_blk0000038e : XORCY
    port map (
      CI => blk00000376_sig000013c1,
      LI => blk00000376_sig000013cd,
      O => blk00000376_sig000013be
    );
  blk00000376_blk0000038d : XORCY
    port map (
      CI => blk00000376_sig0000139b,
      LI => blk00000376_sig000013c2,
      O => blk00000376_sig000013b0
    );
  blk00000376_blk0000038c : MUXCY
    port map (
      CI => blk00000376_sig000013bf,
      DI => blk00000376_sig000013bb,
      S => blk00000376_sig000013cc,
      O => blk00000376_sig000013af
    );
  blk00000376_blk0000038b : XORCY
    port map (
      CI => blk00000376_sig000013bf,
      LI => blk00000376_sig000013cc,
      O => blk00000376_sig000013ae
    );
  blk00000376_blk0000038a : MUXCY
    port map (
      CI => blk00000376_sig000013af,
      DI => blk00000376_sig000013ba,
      S => blk00000376_sig000013cb,
      O => blk00000376_sig000013ad
    );
  blk00000376_blk00000389 : XORCY
    port map (
      CI => blk00000376_sig000013af,
      LI => blk00000376_sig000013cb,
      O => blk00000376_sig000013ac
    );
  blk00000376_blk00000388 : MUXCY
    port map (
      CI => blk00000376_sig000013ad,
      DI => blk00000376_sig000013b9,
      S => blk00000376_sig000013ca,
      O => blk00000376_sig000013ab
    );
  blk00000376_blk00000387 : XORCY
    port map (
      CI => blk00000376_sig000013ad,
      LI => blk00000376_sig000013ca,
      O => blk00000376_sig000013aa
    );
  blk00000376_blk00000386 : MUXCY
    port map (
      CI => blk00000376_sig000013ab,
      DI => blk00000376_sig000013b8,
      S => blk00000376_sig000013c9,
      O => blk00000376_sig000013a9
    );
  blk00000376_blk00000385 : XORCY
    port map (
      CI => blk00000376_sig000013ab,
      LI => blk00000376_sig000013c9,
      O => blk00000376_sig000013a8
    );
  blk00000376_blk00000384 : MUXCY
    port map (
      CI => blk00000376_sig000013a9,
      DI => blk00000376_sig000013b7,
      S => blk00000376_sig000013c8,
      O => blk00000376_sig000013a7
    );
  blk00000376_blk00000383 : XORCY
    port map (
      CI => blk00000376_sig000013a9,
      LI => blk00000376_sig000013c8,
      O => blk00000376_sig000013a6
    );
  blk00000376_blk00000382 : MUXCY
    port map (
      CI => blk00000376_sig000013a7,
      DI => blk00000376_sig000013b6,
      S => blk00000376_sig000013c7,
      O => blk00000376_sig000013a5
    );
  blk00000376_blk00000381 : XORCY
    port map (
      CI => blk00000376_sig000013a7,
      LI => blk00000376_sig000013c7,
      O => blk00000376_sig000013a4
    );
  blk00000376_blk00000380 : MUXCY
    port map (
      CI => blk00000376_sig000013a5,
      DI => blk00000376_sig000013b5,
      S => blk00000376_sig000013c6,
      O => blk00000376_sig000013a3
    );
  blk00000376_blk0000037f : XORCY
    port map (
      CI => blk00000376_sig000013a5,
      LI => blk00000376_sig000013c6,
      O => blk00000376_sig000013a2
    );
  blk00000376_blk0000037e : MUXCY
    port map (
      CI => blk00000376_sig000013a3,
      DI => blk00000376_sig000013b4,
      S => blk00000376_sig000013c5,
      O => blk00000376_sig000013a1
    );
  blk00000376_blk0000037d : XORCY
    port map (
      CI => blk00000376_sig000013a3,
      LI => blk00000376_sig000013c5,
      O => blk00000376_sig000013a0
    );
  blk00000376_blk0000037c : MUXCY
    port map (
      CI => blk00000376_sig000013a1,
      DI => blk00000376_sig000013b3,
      S => blk00000376_sig000013c4,
      O => blk00000376_sig0000139f
    );
  blk00000376_blk0000037b : XORCY
    port map (
      CI => blk00000376_sig000013a1,
      LI => blk00000376_sig000013c4,
      O => blk00000376_sig0000139e
    );
  blk00000376_blk0000037a : MUXCY
    port map (
      CI => blk00000376_sig0000139f,
      DI => blk00000376_sig000013b2,
      S => blk00000376_sig000013c3,
      O => blk00000376_sig0000139d
    );
  blk00000376_blk00000379 : XORCY
    port map (
      CI => blk00000376_sig0000139f,
      LI => blk00000376_sig000013c3,
      O => blk00000376_sig0000139c
    );
  blk00000376_blk00000378 : MUXCY
    port map (
      CI => blk00000376_sig0000139d,
      DI => blk00000376_sig000013b1,
      S => blk00000376_sig000013cf,
      O => blk00000376_sig0000139b
    );
  blk00000376_blk00000377 : XORCY
    port map (
      CI => blk00000376_sig0000139d,
      LI => blk00000376_sig000013cf,
      O => blk00000376_sig0000139a
    );
  blk000003bb_blk000003bc_blk000003bf : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk000003bb_blk000003bc_sig000013e4,
      Q => sig00000111
    );
  blk000003bb_blk000003bc_blk000003be : SRLC32E
    generic map(
      INIT => X"00000000"
    )
    port map (
      CLK => clk,
      D => sig0000027f,
      CE => ce,
      Q => blk000003bb_blk000003bc_sig000013e4,
      Q31 => NLW_blk000003bb_blk000003bc_blk000003be_Q31_UNCONNECTED,
      A(4) => blk000003bb_blk000003bc_sig000013e3,
      A(3) => blk000003bb_blk000003bc_sig000013e3,
      A(2) => blk000003bb_blk000003bc_sig000013e3,
      A(1) => blk000003bb_blk000003bc_sig000013e3,
      A(0) => blk000003bb_blk000003bc_sig000013e3
    );
  blk000003bb_blk000003bc_blk000003bd : VCC
    port map (
      P => blk000003bb_blk000003bc_sig000013e3
    );
  blk000003c0_blk000003c1_blk000003ce : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk000003c0_blk000003c1_sig00001408,
      Q => sig0000010b
    );
  blk000003c0_blk000003c1_blk000003cd : SRLC32E
    generic map(
      INIT => X"00000000"
    )
    port map (
      CLK => clk,
      D => sig0000025f,
      CE => ce,
      Q => blk000003c0_blk000003c1_sig00001408,
      Q31 => NLW_blk000003c0_blk000003c1_blk000003cd_Q31_UNCONNECTED,
      A(4) => blk000003c0_blk000003c1_sig00001402,
      A(3) => blk000003c0_blk000003c1_sig00001402,
      A(2) => blk000003c0_blk000003c1_sig00001402,
      A(1) => blk000003c0_blk000003c1_sig00001402,
      A(0) => blk000003c0_blk000003c1_sig00001402
    );
  blk000003c0_blk000003c1_blk000003cc : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk000003c0_blk000003c1_sig00001407,
      Q => sig0000010a
    );
  blk000003c0_blk000003c1_blk000003cb : SRLC32E
    generic map(
      INIT => X"00000000"
    )
    port map (
      CLK => clk,
      D => sig0000025e,
      CE => ce,
      Q => blk000003c0_blk000003c1_sig00001407,
      Q31 => NLW_blk000003c0_blk000003c1_blk000003cb_Q31_UNCONNECTED,
      A(4) => blk000003c0_blk000003c1_sig00001402,
      A(3) => blk000003c0_blk000003c1_sig00001402,
      A(2) => blk000003c0_blk000003c1_sig00001402,
      A(1) => blk000003c0_blk000003c1_sig00001402,
      A(0) => blk000003c0_blk000003c1_sig00001402
    );
  blk000003c0_blk000003c1_blk000003ca : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk000003c0_blk000003c1_sig00001406,
      Q => sig0000010c
    );
  blk000003c0_blk000003c1_blk000003c9 : SRLC32E
    generic map(
      INIT => X"00000000"
    )
    port map (
      CLK => clk,
      D => sig00000260,
      CE => ce,
      Q => blk000003c0_blk000003c1_sig00001406,
      Q31 => NLW_blk000003c0_blk000003c1_blk000003c9_Q31_UNCONNECTED,
      A(4) => blk000003c0_blk000003c1_sig00001402,
      A(3) => blk000003c0_blk000003c1_sig00001402,
      A(2) => blk000003c0_blk000003c1_sig00001402,
      A(1) => blk000003c0_blk000003c1_sig00001402,
      A(0) => blk000003c0_blk000003c1_sig00001402
    );
  blk000003c0_blk000003c1_blk000003c8 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk000003c0_blk000003c1_sig00001405,
      Q => sig00000108
    );
  blk000003c0_blk000003c1_blk000003c7 : SRLC32E
    generic map(
      INIT => X"00000000"
    )
    port map (
      CLK => clk,
      D => sig0000025c,
      CE => ce,
      Q => blk000003c0_blk000003c1_sig00001405,
      Q31 => NLW_blk000003c0_blk000003c1_blk000003c7_Q31_UNCONNECTED,
      A(4) => blk000003c0_blk000003c1_sig00001402,
      A(3) => blk000003c0_blk000003c1_sig00001402,
      A(2) => blk000003c0_blk000003c1_sig00001402,
      A(1) => blk000003c0_blk000003c1_sig00001402,
      A(0) => blk000003c0_blk000003c1_sig00001402
    );
  blk000003c0_blk000003c1_blk000003c6 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk000003c0_blk000003c1_sig00001404,
      Q => sig00000107
    );
  blk000003c0_blk000003c1_blk000003c5 : SRLC32E
    generic map(
      INIT => X"00000000"
    )
    port map (
      CLK => clk,
      D => sig0000025b,
      CE => ce,
      Q => blk000003c0_blk000003c1_sig00001404,
      Q31 => NLW_blk000003c0_blk000003c1_blk000003c5_Q31_UNCONNECTED,
      A(4) => blk000003c0_blk000003c1_sig00001402,
      A(3) => blk000003c0_blk000003c1_sig00001402,
      A(2) => blk000003c0_blk000003c1_sig00001402,
      A(1) => blk000003c0_blk000003c1_sig00001402,
      A(0) => blk000003c0_blk000003c1_sig00001402
    );
  blk000003c0_blk000003c1_blk000003c4 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk000003c0_blk000003c1_sig00001403,
      Q => sig00000109
    );
  blk000003c0_blk000003c1_blk000003c3 : SRLC32E
    generic map(
      INIT => X"00000000"
    )
    port map (
      CLK => clk,
      D => sig0000025d,
      CE => ce,
      Q => blk000003c0_blk000003c1_sig00001403,
      Q31 => NLW_blk000003c0_blk000003c1_blk000003c3_Q31_UNCONNECTED,
      A(4) => blk000003c0_blk000003c1_sig00001402,
      A(3) => blk000003c0_blk000003c1_sig00001402,
      A(2) => blk000003c0_blk000003c1_sig00001402,
      A(1) => blk000003c0_blk000003c1_sig00001402,
      A(0) => blk000003c0_blk000003c1_sig00001402
    );
  blk000003c0_blk000003c1_blk000003c2 : VCC
    port map (
      P => blk000003c0_blk000003c1_sig00001402
    );
  blk000003cf_blk000003d0_blk000003d4 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk000003cf_blk000003d0_sig00001413,
      Q => sig000001e7
    );
  blk000003cf_blk000003d0_blk000003d3 : SRLC32E
    generic map(
      INIT => X"00000000"
    )
    port map (
      CLK => clk,
      D => sig0000027b,
      CE => ce,
      Q => blk000003cf_blk000003d0_sig00001413,
      Q31 => NLW_blk000003cf_blk000003d0_blk000003d3_Q31_UNCONNECTED,
      A(4) => blk000003cf_blk000003d0_sig00001412,
      A(3) => blk000003cf_blk000003d0_sig00001412,
      A(2) => blk000003cf_blk000003d0_sig00001412,
      A(1) => blk000003cf_blk000003d0_sig00001412,
      A(0) => blk000003cf_blk000003d0_sig00001411
    );
  blk000003cf_blk000003d0_blk000003d2 : VCC
    port map (
      P => blk000003cf_blk000003d0_sig00001412
    );
  blk000003cf_blk000003d0_blk000003d1 : GND
    port map (
      G => blk000003cf_blk000003d0_sig00001411
    );
  blk000003d5_blk000003d6_blk000003da : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk000003d5_blk000003d6_sig0000141f,
      Q => sig00000259
    );
  blk000003d5_blk000003d6_blk000003d9 : SRLC16E
    generic map(
      INIT => X"0000"
    )
    port map (
      A0 => blk000003d5_blk000003d6_sig0000141d,
      A1 => blk000003d5_blk000003d6_sig0000141e,
      A2 => blk000003d5_blk000003d6_sig0000141d,
      A3 => blk000003d5_blk000003d6_sig0000141d,
      CE => ce,
      CLK => clk,
      D => sig0000025a,
      Q => blk000003d5_blk000003d6_sig0000141f,
      Q15 => NLW_blk000003d5_blk000003d6_blk000003d9_Q15_UNCONNECTED
    );
  blk000003d5_blk000003d6_blk000003d8 : VCC
    port map (
      P => blk000003d5_blk000003d6_sig0000141e
    );
  blk000003d5_blk000003d6_blk000003d7 : GND
    port map (
      G => blk000003d5_blk000003d6_sig0000141d
    );
  blk000003db_blk000003dc_blk000003df : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk000003db_blk000003dc_sig00001429,
      Q => sig000000ed
    );
  blk000003db_blk000003dc_blk000003de : SRLC32E
    generic map(
      INIT => X"00000000"
    )
    port map (
      CLK => clk,
      D => sig000001eb,
      CE => ce,
      Q => blk000003db_blk000003dc_sig00001429,
      Q31 => NLW_blk000003db_blk000003dc_blk000003de_Q31_UNCONNECTED,
      A(4) => blk000003db_blk000003dc_sig00001428,
      A(3) => blk000003db_blk000003dc_sig00001428,
      A(2) => blk000003db_blk000003dc_sig00001428,
      A(1) => blk000003db_blk000003dc_sig00001428,
      A(0) => blk000003db_blk000003dc_sig00001428
    );
  blk000003db_blk000003dc_blk000003dd : VCC
    port map (
      P => blk000003db_blk000003dc_sig00001428
    );
  blk000003e0_blk000003e1_blk000003e7 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk000003e0_blk000003e1_sig00001439,
      Q => sig00000252
    );
  blk000003e0_blk000003e1_blk000003e6 : SRLC32E
    generic map(
      INIT => X"00000000"
    )
    port map (
      CLK => clk,
      D => sig00000254,
      CE => ce,
      Q => blk000003e0_blk000003e1_sig00001439,
      Q31 => NLW_blk000003e0_blk000003e1_blk000003e6_Q31_UNCONNECTED,
      A(4) => blk000003e0_blk000003e1_sig00001437,
      A(3) => blk000003e0_blk000003e1_sig00001437,
      A(2) => blk000003e0_blk000003e1_sig00001437,
      A(1) => blk000003e0_blk000003e1_sig00001437,
      A(0) => blk000003e0_blk000003e1_sig00001436
    );
  blk000003e0_blk000003e1_blk000003e5 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk000003e0_blk000003e1_sig00001438,
      Q => sig00000251
    );
  blk000003e0_blk000003e1_blk000003e4 : SRLC32E
    generic map(
      INIT => X"00000000"
    )
    port map (
      CLK => clk,
      D => sig00000253,
      CE => ce,
      Q => blk000003e0_blk000003e1_sig00001438,
      Q31 => NLW_blk000003e0_blk000003e1_blk000003e4_Q31_UNCONNECTED,
      A(4) => blk000003e0_blk000003e1_sig00001437,
      A(3) => blk000003e0_blk000003e1_sig00001437,
      A(2) => blk000003e0_blk000003e1_sig00001437,
      A(1) => blk000003e0_blk000003e1_sig00001437,
      A(0) => blk000003e0_blk000003e1_sig00001436
    );
  blk000003e0_blk000003e1_blk000003e3 : VCC
    port map (
      P => blk000003e0_blk000003e1_sig00001437
    );
  blk000003e0_blk000003e1_blk000003e2 : GND
    port map (
      G => blk000003e0_blk000003e1_sig00001436
    );
  blk000003e8_blk000003e9_blk000003f2 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk000003e8_blk000003e9_sig00001452,
      Q => sig00000110
    );
  blk000003e8_blk000003e9_blk000003f1 : SRLC32E
    generic map(
      INIT => X"00000000"
    )
    port map (
      CLK => clk,
      D => sig00000258,
      CE => ce,
      Q => blk000003e8_blk000003e9_sig00001452,
      Q31 => NLW_blk000003e8_blk000003e9_blk000003f1_Q31_UNCONNECTED,
      A(4) => blk000003e8_blk000003e9_sig0000144e,
      A(3) => blk000003e8_blk000003e9_sig0000144e,
      A(2) => blk000003e8_blk000003e9_sig0000144e,
      A(1) => blk000003e8_blk000003e9_sig0000144e,
      A(0) => blk000003e8_blk000003e9_sig0000144e
    );
  blk000003e8_blk000003e9_blk000003f0 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk000003e8_blk000003e9_sig00001451,
      Q => sig0000010f
    );
  blk000003e8_blk000003e9_blk000003ef : SRLC32E
    generic map(
      INIT => X"00000000"
    )
    port map (
      CLK => clk,
      D => sig00000257,
      CE => ce,
      Q => blk000003e8_blk000003e9_sig00001451,
      Q31 => NLW_blk000003e8_blk000003e9_blk000003ef_Q31_UNCONNECTED,
      A(4) => blk000003e8_blk000003e9_sig0000144e,
      A(3) => blk000003e8_blk000003e9_sig0000144e,
      A(2) => blk000003e8_blk000003e9_sig0000144e,
      A(1) => blk000003e8_blk000003e9_sig0000144e,
      A(0) => blk000003e8_blk000003e9_sig0000144e
    );
  blk000003e8_blk000003e9_blk000003ee : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk000003e8_blk000003e9_sig00001450,
      Q => sig0000010e
    );
  blk000003e8_blk000003e9_blk000003ed : SRLC32E
    generic map(
      INIT => X"00000000"
    )
    port map (
      CLK => clk,
      D => sig00000256,
      CE => ce,
      Q => blk000003e8_blk000003e9_sig00001450,
      Q31 => NLW_blk000003e8_blk000003e9_blk000003ed_Q31_UNCONNECTED,
      A(4) => blk000003e8_blk000003e9_sig0000144e,
      A(3) => blk000003e8_blk000003e9_sig0000144e,
      A(2) => blk000003e8_blk000003e9_sig0000144e,
      A(1) => blk000003e8_blk000003e9_sig0000144e,
      A(0) => blk000003e8_blk000003e9_sig0000144e
    );
  blk000003e8_blk000003e9_blk000003ec : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk000003e8_blk000003e9_sig0000144f,
      Q => sig0000010d
    );
  blk000003e8_blk000003e9_blk000003eb : SRLC32E
    generic map(
      INIT => X"00000000"
    )
    port map (
      CLK => clk,
      D => sig00000255,
      CE => ce,
      Q => blk000003e8_blk000003e9_sig0000144f,
      Q31 => NLW_blk000003e8_blk000003e9_blk000003eb_Q31_UNCONNECTED,
      A(4) => blk000003e8_blk000003e9_sig0000144e,
      A(3) => blk000003e8_blk000003e9_sig0000144e,
      A(2) => blk000003e8_blk000003e9_sig0000144e,
      A(1) => blk000003e8_blk000003e9_sig0000144e,
      A(0) => blk000003e8_blk000003e9_sig0000144e
    );
  blk000003e8_blk000003e9_blk000003ea : VCC
    port map (
      P => blk000003e8_blk000003e9_sig0000144e
    );
  blk000004a0_blk000004a1_blk000004a4 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk000004a0_blk000004a1_sig00001463,
      Q => sig00000491
    );
  blk000004a0_blk000004a1_blk000004a3 : SRLC16E
    generic map(
      INIT => X"0000"
    )
    port map (
      A0 => blk000004a0_blk000004a1_sig00001462,
      A1 => blk000004a0_blk000004a1_sig00001462,
      A2 => blk000004a0_blk000004a1_sig00001462,
      A3 => blk000004a0_blk000004a1_sig00001462,
      CE => ce,
      CLK => clk,
      D => sig00000492,
      Q => blk000004a0_blk000004a1_sig00001463,
      Q15 => NLW_blk000004a0_blk000004a1_blk000004a3_Q15_UNCONNECTED
    );
  blk000004a0_blk000004a1_blk000004a2 : GND
    port map (
      G => blk000004a0_blk000004a1_sig00001462
    );
  blk000004a5_blk000004a6_blk000004a9 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk000004a5_blk000004a6_sig00001474,
      Q => sig00000490
    );
  blk000004a5_blk000004a6_blk000004a8 : SRLC16E
    generic map(
      INIT => X"0000"
    )
    port map (
      A0 => blk000004a5_blk000004a6_sig00001473,
      A1 => blk000004a5_blk000004a6_sig00001473,
      A2 => blk000004a5_blk000004a6_sig00001473,
      A3 => blk000004a5_blk000004a6_sig00001473,
      CE => ce,
      CLK => clk,
      D => sig00000491,
      Q => blk000004a5_blk000004a6_sig00001474,
      Q15 => NLW_blk000004a5_blk000004a6_blk000004a8_Q15_UNCONNECTED
    );
  blk000004a5_blk000004a6_blk000004a7 : GND
    port map (
      G => blk000004a5_blk000004a6_sig00001473
    );
  blk000004aa_blk000004ab_blk000004ae : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk000004aa_blk000004ab_sig00001485,
      Q => sig00000001
    );
  blk000004aa_blk000004ab_blk000004ad : SRLC16E
    generic map(
      INIT => X"0000"
    )
    port map (
      A0 => blk000004aa_blk000004ab_sig00001484,
      A1 => blk000004aa_blk000004ab_sig00001484,
      A2 => blk000004aa_blk000004ab_sig00001484,
      A3 => blk000004aa_blk000004ab_sig00001484,
      CE => ce,
      CLK => clk,
      D => sig000000a3,
      Q => blk000004aa_blk000004ab_sig00001485,
      Q15 => NLW_blk000004aa_blk000004ab_blk000004ad_Q15_UNCONNECTED
    );
  blk000004aa_blk000004ab_blk000004ac : GND
    port map (
      G => blk000004aa_blk000004ab_sig00001484
    );
  blk000004af_blk000004b0_blk000004b3 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk000004af_blk000004b0_sig00001496,
      Q => sig000000a1
    );
  blk000004af_blk000004b0_blk000004b2 : SRLC16E
    generic map(
      INIT => X"0000"
    )
    port map (
      A0 => blk000004af_blk000004b0_sig00001495,
      A1 => blk000004af_blk000004b0_sig00001495,
      A2 => blk000004af_blk000004b0_sig00001495,
      A3 => blk000004af_blk000004b0_sig00001495,
      CE => ce,
      CLK => clk,
      D => sig00000115,
      Q => blk000004af_blk000004b0_sig00001496,
      Q15 => NLW_blk000004af_blk000004b0_blk000004b2_Q15_UNCONNECTED
    );
  blk000004af_blk000004b0_blk000004b1 : GND
    port map (
      G => blk000004af_blk000004b0_sig00001495
    );
  blk000004b4_blk000004b5_blk000004b9 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk000004b4_blk000004b5_sig000014a2,
      Q => sig0000048f
    );
  blk000004b4_blk000004b5_blk000004b8 : SRLC16E
    generic map(
      INIT => X"0000"
    )
    port map (
      A0 => blk000004b4_blk000004b5_sig000014a0,
      A1 => blk000004b4_blk000004b5_sig000014a1,
      A2 => blk000004b4_blk000004b5_sig000014a1,
      A3 => blk000004b4_blk000004b5_sig000014a1,
      CE => ce,
      CLK => clk,
      D => sig00000490,
      Q => blk000004b4_blk000004b5_sig000014a2,
      Q15 => NLW_blk000004b4_blk000004b5_blk000004b8_Q15_UNCONNECTED
    );
  blk000004b4_blk000004b5_blk000004b7 : VCC
    port map (
      P => blk000004b4_blk000004b5_sig000014a1
    );
  blk000004b4_blk000004b5_blk000004b6 : GND
    port map (
      G => blk000004b4_blk000004b5_sig000014a0
    );
  blk000004ba_blk000004bb_blk000004d9 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk000004ba_blk000004bb_sig000014ef,
      Q => sig00000470
    );
  blk000004ba_blk000004bb_blk000004d8 : SRLC16E
    generic map(
      INIT => X"0000"
    )
    port map (
      A0 => blk000004ba_blk000004bb_sig000014e0,
      A1 => blk000004ba_blk000004bb_sig000014e1,
      A2 => blk000004ba_blk000004bb_sig000014e1,
      A3 => blk000004ba_blk000004bb_sig000014e1,
      CE => ce,
      CLK => clk,
      D => sig00000454,
      Q => blk000004ba_blk000004bb_sig000014ef,
      Q15 => NLW_blk000004ba_blk000004bb_blk000004d8_Q15_UNCONNECTED
    );
  blk000004ba_blk000004bb_blk000004d7 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk000004ba_blk000004bb_sig000014ee,
      Q => sig0000046f
    );
  blk000004ba_blk000004bb_blk000004d6 : SRLC16E
    generic map(
      INIT => X"0000"
    )
    port map (
      A0 => blk000004ba_blk000004bb_sig000014e0,
      A1 => blk000004ba_blk000004bb_sig000014e1,
      A2 => blk000004ba_blk000004bb_sig000014e1,
      A3 => blk000004ba_blk000004bb_sig000014e1,
      CE => ce,
      CLK => clk,
      D => sig00000453,
      Q => blk000004ba_blk000004bb_sig000014ee,
      Q15 => NLW_blk000004ba_blk000004bb_blk000004d6_Q15_UNCONNECTED
    );
  blk000004ba_blk000004bb_blk000004d5 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk000004ba_blk000004bb_sig000014ed,
      Q => sig00000471
    );
  blk000004ba_blk000004bb_blk000004d4 : SRLC16E
    generic map(
      INIT => X"0000"
    )
    port map (
      A0 => blk000004ba_blk000004bb_sig000014e0,
      A1 => blk000004ba_blk000004bb_sig000014e1,
      A2 => blk000004ba_blk000004bb_sig000014e1,
      A3 => blk000004ba_blk000004bb_sig000014e1,
      CE => ce,
      CLK => clk,
      D => sig00000455,
      Q => blk000004ba_blk000004bb_sig000014ed,
      Q15 => NLW_blk000004ba_blk000004bb_blk000004d4_Q15_UNCONNECTED
    );
  blk000004ba_blk000004bb_blk000004d3 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk000004ba_blk000004bb_sig000014ec,
      Q => sig0000046e
    );
  blk000004ba_blk000004bb_blk000004d2 : SRLC16E
    generic map(
      INIT => X"0000"
    )
    port map (
      A0 => blk000004ba_blk000004bb_sig000014e0,
      A1 => blk000004ba_blk000004bb_sig000014e1,
      A2 => blk000004ba_blk000004bb_sig000014e1,
      A3 => blk000004ba_blk000004bb_sig000014e1,
      CE => ce,
      CLK => clk,
      D => sig00000452,
      Q => blk000004ba_blk000004bb_sig000014ec,
      Q15 => NLW_blk000004ba_blk000004bb_blk000004d2_Q15_UNCONNECTED
    );
  blk000004ba_blk000004bb_blk000004d1 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk000004ba_blk000004bb_sig000014eb,
      Q => sig0000046d
    );
  blk000004ba_blk000004bb_blk000004d0 : SRLC16E
    generic map(
      INIT => X"0000"
    )
    port map (
      A0 => blk000004ba_blk000004bb_sig000014e0,
      A1 => blk000004ba_blk000004bb_sig000014e1,
      A2 => blk000004ba_blk000004bb_sig000014e1,
      A3 => blk000004ba_blk000004bb_sig000014e1,
      CE => ce,
      CLK => clk,
      D => sig00000451,
      Q => blk000004ba_blk000004bb_sig000014eb,
      Q15 => NLW_blk000004ba_blk000004bb_blk000004d0_Q15_UNCONNECTED
    );
  blk000004ba_blk000004bb_blk000004cf : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk000004ba_blk000004bb_sig000014ea,
      Q => sig0000046c
    );
  blk000004ba_blk000004bb_blk000004ce : SRLC16E
    generic map(
      INIT => X"0000"
    )
    port map (
      A0 => blk000004ba_blk000004bb_sig000014e0,
      A1 => blk000004ba_blk000004bb_sig000014e1,
      A2 => blk000004ba_blk000004bb_sig000014e1,
      A3 => blk000004ba_blk000004bb_sig000014e1,
      CE => ce,
      CLK => clk,
      D => sig00000450,
      Q => blk000004ba_blk000004bb_sig000014ea,
      Q15 => NLW_blk000004ba_blk000004bb_blk000004ce_Q15_UNCONNECTED
    );
  blk000004ba_blk000004bb_blk000004cd : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk000004ba_blk000004bb_sig000014e9,
      Q => sig0000046b
    );
  blk000004ba_blk000004bb_blk000004cc : SRLC16E
    generic map(
      INIT => X"0000"
    )
    port map (
      A0 => blk000004ba_blk000004bb_sig000014e0,
      A1 => blk000004ba_blk000004bb_sig000014e1,
      A2 => blk000004ba_blk000004bb_sig000014e1,
      A3 => blk000004ba_blk000004bb_sig000014e1,
      CE => ce,
      CLK => clk,
      D => sig0000044f,
      Q => blk000004ba_blk000004bb_sig000014e9,
      Q15 => NLW_blk000004ba_blk000004bb_blk000004cc_Q15_UNCONNECTED
    );
  blk000004ba_blk000004bb_blk000004cb : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk000004ba_blk000004bb_sig000014e8,
      Q => sig00000469
    );
  blk000004ba_blk000004bb_blk000004ca : SRLC16E
    generic map(
      INIT => X"0000"
    )
    port map (
      A0 => blk000004ba_blk000004bb_sig000014e0,
      A1 => blk000004ba_blk000004bb_sig000014e1,
      A2 => blk000004ba_blk000004bb_sig000014e1,
      A3 => blk000004ba_blk000004bb_sig000014e1,
      CE => ce,
      CLK => clk,
      D => sig0000044d,
      Q => blk000004ba_blk000004bb_sig000014e8,
      Q15 => NLW_blk000004ba_blk000004bb_blk000004ca_Q15_UNCONNECTED
    );
  blk000004ba_blk000004bb_blk000004c9 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk000004ba_blk000004bb_sig000014e7,
      Q => sig00000468
    );
  blk000004ba_blk000004bb_blk000004c8 : SRLC16E
    generic map(
      INIT => X"0000"
    )
    port map (
      A0 => blk000004ba_blk000004bb_sig000014e0,
      A1 => blk000004ba_blk000004bb_sig000014e1,
      A2 => blk000004ba_blk000004bb_sig000014e1,
      A3 => blk000004ba_blk000004bb_sig000014e1,
      CE => ce,
      CLK => clk,
      D => sig0000044c,
      Q => blk000004ba_blk000004bb_sig000014e7,
      Q15 => NLW_blk000004ba_blk000004bb_blk000004c8_Q15_UNCONNECTED
    );
  blk000004ba_blk000004bb_blk000004c7 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk000004ba_blk000004bb_sig000014e6,
      Q => sig0000046a
    );
  blk000004ba_blk000004bb_blk000004c6 : SRLC16E
    generic map(
      INIT => X"0000"
    )
    port map (
      A0 => blk000004ba_blk000004bb_sig000014e0,
      A1 => blk000004ba_blk000004bb_sig000014e1,
      A2 => blk000004ba_blk000004bb_sig000014e1,
      A3 => blk000004ba_blk000004bb_sig000014e1,
      CE => ce,
      CLK => clk,
      D => sig0000044e,
      Q => blk000004ba_blk000004bb_sig000014e6,
      Q15 => NLW_blk000004ba_blk000004bb_blk000004c6_Q15_UNCONNECTED
    );
  blk000004ba_blk000004bb_blk000004c5 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk000004ba_blk000004bb_sig000014e5,
      Q => sig00000467
    );
  blk000004ba_blk000004bb_blk000004c4 : SRLC16E
    generic map(
      INIT => X"0000"
    )
    port map (
      A0 => blk000004ba_blk000004bb_sig000014e0,
      A1 => blk000004ba_blk000004bb_sig000014e1,
      A2 => blk000004ba_blk000004bb_sig000014e1,
      A3 => blk000004ba_blk000004bb_sig000014e1,
      CE => ce,
      CLK => clk,
      D => sig0000044b,
      Q => blk000004ba_blk000004bb_sig000014e5,
      Q15 => NLW_blk000004ba_blk000004bb_blk000004c4_Q15_UNCONNECTED
    );
  blk000004ba_blk000004bb_blk000004c3 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk000004ba_blk000004bb_sig000014e4,
      Q => sig00000466
    );
  blk000004ba_blk000004bb_blk000004c2 : SRLC16E
    generic map(
      INIT => X"0000"
    )
    port map (
      A0 => blk000004ba_blk000004bb_sig000014e0,
      A1 => blk000004ba_blk000004bb_sig000014e1,
      A2 => blk000004ba_blk000004bb_sig000014e1,
      A3 => blk000004ba_blk000004bb_sig000014e1,
      CE => ce,
      CLK => clk,
      D => sig0000044a,
      Q => blk000004ba_blk000004bb_sig000014e4,
      Q15 => NLW_blk000004ba_blk000004bb_blk000004c2_Q15_UNCONNECTED
    );
  blk000004ba_blk000004bb_blk000004c1 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk000004ba_blk000004bb_sig000014e3,
      Q => sig00000465
    );
  blk000004ba_blk000004bb_blk000004c0 : SRLC16E
    generic map(
      INIT => X"0000"
    )
    port map (
      A0 => blk000004ba_blk000004bb_sig000014e0,
      A1 => blk000004ba_blk000004bb_sig000014e1,
      A2 => blk000004ba_blk000004bb_sig000014e1,
      A3 => blk000004ba_blk000004bb_sig000014e1,
      CE => ce,
      CLK => clk,
      D => sig00000449,
      Q => blk000004ba_blk000004bb_sig000014e3,
      Q15 => NLW_blk000004ba_blk000004bb_blk000004c0_Q15_UNCONNECTED
    );
  blk000004ba_blk000004bb_blk000004bf : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk000004ba_blk000004bb_sig000014e2,
      Q => sig00000464
    );
  blk000004ba_blk000004bb_blk000004be : SRLC16E
    generic map(
      INIT => X"0000"
    )
    port map (
      A0 => blk000004ba_blk000004bb_sig000014e0,
      A1 => blk000004ba_blk000004bb_sig000014e1,
      A2 => blk000004ba_blk000004bb_sig000014e1,
      A3 => blk000004ba_blk000004bb_sig000014e1,
      CE => ce,
      CLK => clk,
      D => sig00000448,
      Q => blk000004ba_blk000004bb_sig000014e2,
      Q15 => NLW_blk000004ba_blk000004bb_blk000004be_Q15_UNCONNECTED
    );
  blk000004ba_blk000004bb_blk000004bd : VCC
    port map (
      P => blk000004ba_blk000004bb_sig000014e1
    );
  blk000004ba_blk000004bb_blk000004bc : GND
    port map (
      G => blk000004ba_blk000004bb_sig000014e0
    );
  blk000004da_blk000004db_blk000004f9 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk000004da_blk000004db_sig0000153c,
      Q => sig00000462
    );
  blk000004da_blk000004db_blk000004f8 : SRLC16E
    generic map(
      INIT => X"0000"
    )
    port map (
      A0 => blk000004da_blk000004db_sig0000152d,
      A1 => blk000004da_blk000004db_sig0000152e,
      A2 => blk000004da_blk000004db_sig0000152e,
      A3 => blk000004da_blk000004db_sig0000152e,
      CE => ce,
      CLK => clk,
      D => sig00000400,
      Q => blk000004da_blk000004db_sig0000153c,
      Q15 => NLW_blk000004da_blk000004db_blk000004f8_Q15_UNCONNECTED
    );
  blk000004da_blk000004db_blk000004f7 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk000004da_blk000004db_sig0000153b,
      Q => sig00000461
    );
  blk000004da_blk000004db_blk000004f6 : SRLC16E
    generic map(
      INIT => X"0000"
    )
    port map (
      A0 => blk000004da_blk000004db_sig0000152d,
      A1 => blk000004da_blk000004db_sig0000152e,
      A2 => blk000004da_blk000004db_sig0000152e,
      A3 => blk000004da_blk000004db_sig0000152e,
      CE => ce,
      CLK => clk,
      D => sig000003ff,
      Q => blk000004da_blk000004db_sig0000153b,
      Q15 => NLW_blk000004da_blk000004db_blk000004f6_Q15_UNCONNECTED
    );
  blk000004da_blk000004db_blk000004f5 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk000004da_blk000004db_sig0000153a,
      Q => sig00000463
    );
  blk000004da_blk000004db_blk000004f4 : SRLC16E
    generic map(
      INIT => X"0000"
    )
    port map (
      A0 => blk000004da_blk000004db_sig0000152d,
      A1 => blk000004da_blk000004db_sig0000152e,
      A2 => blk000004da_blk000004db_sig0000152e,
      A3 => blk000004da_blk000004db_sig0000152e,
      CE => ce,
      CLK => clk,
      D => sig00000401,
      Q => blk000004da_blk000004db_sig0000153a,
      Q15 => NLW_blk000004da_blk000004db_blk000004f4_Q15_UNCONNECTED
    );
  blk000004da_blk000004db_blk000004f3 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk000004da_blk000004db_sig00001539,
      Q => sig00000460
    );
  blk000004da_blk000004db_blk000004f2 : SRLC16E
    generic map(
      INIT => X"0000"
    )
    port map (
      A0 => blk000004da_blk000004db_sig0000152d,
      A1 => blk000004da_blk000004db_sig0000152e,
      A2 => blk000004da_blk000004db_sig0000152e,
      A3 => blk000004da_blk000004db_sig0000152e,
      CE => ce,
      CLK => clk,
      D => sig000003fe,
      Q => blk000004da_blk000004db_sig00001539,
      Q15 => NLW_blk000004da_blk000004db_blk000004f2_Q15_UNCONNECTED
    );
  blk000004da_blk000004db_blk000004f1 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk000004da_blk000004db_sig00001538,
      Q => sig0000045f
    );
  blk000004da_blk000004db_blk000004f0 : SRLC16E
    generic map(
      INIT => X"0000"
    )
    port map (
      A0 => blk000004da_blk000004db_sig0000152d,
      A1 => blk000004da_blk000004db_sig0000152e,
      A2 => blk000004da_blk000004db_sig0000152e,
      A3 => blk000004da_blk000004db_sig0000152e,
      CE => ce,
      CLK => clk,
      D => sig000003fd,
      Q => blk000004da_blk000004db_sig00001538,
      Q15 => NLW_blk000004da_blk000004db_blk000004f0_Q15_UNCONNECTED
    );
  blk000004da_blk000004db_blk000004ef : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk000004da_blk000004db_sig00001537,
      Q => sig0000045e
    );
  blk000004da_blk000004db_blk000004ee : SRLC16E
    generic map(
      INIT => X"0000"
    )
    port map (
      A0 => blk000004da_blk000004db_sig0000152d,
      A1 => blk000004da_blk000004db_sig0000152e,
      A2 => blk000004da_blk000004db_sig0000152e,
      A3 => blk000004da_blk000004db_sig0000152e,
      CE => ce,
      CLK => clk,
      D => sig000003fc,
      Q => blk000004da_blk000004db_sig00001537,
      Q15 => NLW_blk000004da_blk000004db_blk000004ee_Q15_UNCONNECTED
    );
  blk000004da_blk000004db_blk000004ed : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk000004da_blk000004db_sig00001536,
      Q => sig0000045d
    );
  blk000004da_blk000004db_blk000004ec : SRLC16E
    generic map(
      INIT => X"0000"
    )
    port map (
      A0 => blk000004da_blk000004db_sig0000152d,
      A1 => blk000004da_blk000004db_sig0000152e,
      A2 => blk000004da_blk000004db_sig0000152e,
      A3 => blk000004da_blk000004db_sig0000152e,
      CE => ce,
      CLK => clk,
      D => sig000003fb,
      Q => blk000004da_blk000004db_sig00001536,
      Q15 => NLW_blk000004da_blk000004db_blk000004ec_Q15_UNCONNECTED
    );
  blk000004da_blk000004db_blk000004eb : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk000004da_blk000004db_sig00001535,
      Q => sig0000045b
    );
  blk000004da_blk000004db_blk000004ea : SRLC16E
    generic map(
      INIT => X"0000"
    )
    port map (
      A0 => blk000004da_blk000004db_sig0000152d,
      A1 => blk000004da_blk000004db_sig0000152e,
      A2 => blk000004da_blk000004db_sig0000152e,
      A3 => blk000004da_blk000004db_sig0000152e,
      CE => ce,
      CLK => clk,
      D => sig000003f9,
      Q => blk000004da_blk000004db_sig00001535,
      Q15 => NLW_blk000004da_blk000004db_blk000004ea_Q15_UNCONNECTED
    );
  blk000004da_blk000004db_blk000004e9 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk000004da_blk000004db_sig00001534,
      Q => sig0000045a
    );
  blk000004da_blk000004db_blk000004e8 : SRLC16E
    generic map(
      INIT => X"0000"
    )
    port map (
      A0 => blk000004da_blk000004db_sig0000152d,
      A1 => blk000004da_blk000004db_sig0000152e,
      A2 => blk000004da_blk000004db_sig0000152e,
      A3 => blk000004da_blk000004db_sig0000152e,
      CE => ce,
      CLK => clk,
      D => sig000003f8,
      Q => blk000004da_blk000004db_sig00001534,
      Q15 => NLW_blk000004da_blk000004db_blk000004e8_Q15_UNCONNECTED
    );
  blk000004da_blk000004db_blk000004e7 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk000004da_blk000004db_sig00001533,
      Q => sig0000045c
    );
  blk000004da_blk000004db_blk000004e6 : SRLC16E
    generic map(
      INIT => X"0000"
    )
    port map (
      A0 => blk000004da_blk000004db_sig0000152d,
      A1 => blk000004da_blk000004db_sig0000152e,
      A2 => blk000004da_blk000004db_sig0000152e,
      A3 => blk000004da_blk000004db_sig0000152e,
      CE => ce,
      CLK => clk,
      D => sig000003fa,
      Q => blk000004da_blk000004db_sig00001533,
      Q15 => NLW_blk000004da_blk000004db_blk000004e6_Q15_UNCONNECTED
    );
  blk000004da_blk000004db_blk000004e5 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk000004da_blk000004db_sig00001532,
      Q => sig00000459
    );
  blk000004da_blk000004db_blk000004e4 : SRLC16E
    generic map(
      INIT => X"0000"
    )
    port map (
      A0 => blk000004da_blk000004db_sig0000152d,
      A1 => blk000004da_blk000004db_sig0000152e,
      A2 => blk000004da_blk000004db_sig0000152e,
      A3 => blk000004da_blk000004db_sig0000152e,
      CE => ce,
      CLK => clk,
      D => sig000003f7,
      Q => blk000004da_blk000004db_sig00001532,
      Q15 => NLW_blk000004da_blk000004db_blk000004e4_Q15_UNCONNECTED
    );
  blk000004da_blk000004db_blk000004e3 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk000004da_blk000004db_sig00001531,
      Q => sig00000458
    );
  blk000004da_blk000004db_blk000004e2 : SRLC16E
    generic map(
      INIT => X"0000"
    )
    port map (
      A0 => blk000004da_blk000004db_sig0000152d,
      A1 => blk000004da_blk000004db_sig0000152e,
      A2 => blk000004da_blk000004db_sig0000152e,
      A3 => blk000004da_blk000004db_sig0000152e,
      CE => ce,
      CLK => clk,
      D => sig000003f6,
      Q => blk000004da_blk000004db_sig00001531,
      Q15 => NLW_blk000004da_blk000004db_blk000004e2_Q15_UNCONNECTED
    );
  blk000004da_blk000004db_blk000004e1 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk000004da_blk000004db_sig00001530,
      Q => sig00000457
    );
  blk000004da_blk000004db_blk000004e0 : SRLC16E
    generic map(
      INIT => X"0000"
    )
    port map (
      A0 => blk000004da_blk000004db_sig0000152d,
      A1 => blk000004da_blk000004db_sig0000152e,
      A2 => blk000004da_blk000004db_sig0000152e,
      A3 => blk000004da_blk000004db_sig0000152e,
      CE => ce,
      CLK => clk,
      D => sig000003f5,
      Q => blk000004da_blk000004db_sig00001530,
      Q15 => NLW_blk000004da_blk000004db_blk000004e0_Q15_UNCONNECTED
    );
  blk000004da_blk000004db_blk000004df : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk000004da_blk000004db_sig0000152f,
      Q => sig00000456
    );
  blk000004da_blk000004db_blk000004de : SRLC16E
    generic map(
      INIT => X"0000"
    )
    port map (
      A0 => blk000004da_blk000004db_sig0000152d,
      A1 => blk000004da_blk000004db_sig0000152e,
      A2 => blk000004da_blk000004db_sig0000152e,
      A3 => blk000004da_blk000004db_sig0000152e,
      CE => ce,
      CLK => clk,
      D => sig000003f4,
      Q => blk000004da_blk000004db_sig0000152f,
      Q15 => NLW_blk000004da_blk000004db_blk000004de_Q15_UNCONNECTED
    );
  blk000004da_blk000004db_blk000004dd : VCC
    port map (
      P => blk000004da_blk000004db_sig0000152e
    );
  blk000004da_blk000004db_blk000004dc : GND
    port map (
      G => blk000004da_blk000004db_sig0000152d
    );
  blk000004fa_blk000004fb_blk00000519 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk000004fa_blk000004fb_sig00001589,
      Q => sig0000041c
    );
  blk000004fa_blk000004fb_blk00000518 : SRLC16E
    generic map(
      INIT => X"0000"
    )
    port map (
      A0 => blk000004fa_blk000004fb_sig0000157a,
      A1 => blk000004fa_blk000004fb_sig0000157b,
      A2 => blk000004fa_blk000004fb_sig0000157b,
      A3 => blk000004fa_blk000004fb_sig0000157b,
      CE => ce,
      CLK => clk,
      D => sig0000042a,
      Q => blk000004fa_blk000004fb_sig00001589,
      Q15 => NLW_blk000004fa_blk000004fb_blk00000518_Q15_UNCONNECTED
    );
  blk000004fa_blk000004fb_blk00000517 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk000004fa_blk000004fb_sig00001588,
      Q => sig0000041b
    );
  blk000004fa_blk000004fb_blk00000516 : SRLC16E
    generic map(
      INIT => X"0000"
    )
    port map (
      A0 => blk000004fa_blk000004fb_sig0000157a,
      A1 => blk000004fa_blk000004fb_sig0000157b,
      A2 => blk000004fa_blk000004fb_sig0000157b,
      A3 => blk000004fa_blk000004fb_sig0000157b,
      CE => ce,
      CLK => clk,
      D => sig00000429,
      Q => blk000004fa_blk000004fb_sig00001588,
      Q15 => NLW_blk000004fa_blk000004fb_blk00000516_Q15_UNCONNECTED
    );
  blk000004fa_blk000004fb_blk00000515 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk000004fa_blk000004fb_sig00001587,
      Q => sig0000041d
    );
  blk000004fa_blk000004fb_blk00000514 : SRLC16E
    generic map(
      INIT => X"0000"
    )
    port map (
      A0 => blk000004fa_blk000004fb_sig0000157a,
      A1 => blk000004fa_blk000004fb_sig0000157b,
      A2 => blk000004fa_blk000004fb_sig0000157b,
      A3 => blk000004fa_blk000004fb_sig0000157b,
      CE => ce,
      CLK => clk,
      D => sig0000042b,
      Q => blk000004fa_blk000004fb_sig00001587,
      Q15 => NLW_blk000004fa_blk000004fb_blk00000514_Q15_UNCONNECTED
    );
  blk000004fa_blk000004fb_blk00000513 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk000004fa_blk000004fb_sig00001586,
      Q => sig0000041a
    );
  blk000004fa_blk000004fb_blk00000512 : SRLC16E
    generic map(
      INIT => X"0000"
    )
    port map (
      A0 => blk000004fa_blk000004fb_sig0000157a,
      A1 => blk000004fa_blk000004fb_sig0000157b,
      A2 => blk000004fa_blk000004fb_sig0000157b,
      A3 => blk000004fa_blk000004fb_sig0000157b,
      CE => ce,
      CLK => clk,
      D => sig00000428,
      Q => blk000004fa_blk000004fb_sig00001586,
      Q15 => NLW_blk000004fa_blk000004fb_blk00000512_Q15_UNCONNECTED
    );
  blk000004fa_blk000004fb_blk00000511 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk000004fa_blk000004fb_sig00001585,
      Q => sig00000419
    );
  blk000004fa_blk000004fb_blk00000510 : SRLC16E
    generic map(
      INIT => X"0000"
    )
    port map (
      A0 => blk000004fa_blk000004fb_sig0000157a,
      A1 => blk000004fa_blk000004fb_sig0000157b,
      A2 => blk000004fa_blk000004fb_sig0000157b,
      A3 => blk000004fa_blk000004fb_sig0000157b,
      CE => ce,
      CLK => clk,
      D => sig00000427,
      Q => blk000004fa_blk000004fb_sig00001585,
      Q15 => NLW_blk000004fa_blk000004fb_blk00000510_Q15_UNCONNECTED
    );
  blk000004fa_blk000004fb_blk0000050f : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk000004fa_blk000004fb_sig00001584,
      Q => sig00000418
    );
  blk000004fa_blk000004fb_blk0000050e : SRLC16E
    generic map(
      INIT => X"0000"
    )
    port map (
      A0 => blk000004fa_blk000004fb_sig0000157a,
      A1 => blk000004fa_blk000004fb_sig0000157b,
      A2 => blk000004fa_blk000004fb_sig0000157b,
      A3 => blk000004fa_blk000004fb_sig0000157b,
      CE => ce,
      CLK => clk,
      D => sig00000426,
      Q => blk000004fa_blk000004fb_sig00001584,
      Q15 => NLW_blk000004fa_blk000004fb_blk0000050e_Q15_UNCONNECTED
    );
  blk000004fa_blk000004fb_blk0000050d : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk000004fa_blk000004fb_sig00001583,
      Q => sig00000417
    );
  blk000004fa_blk000004fb_blk0000050c : SRLC16E
    generic map(
      INIT => X"0000"
    )
    port map (
      A0 => blk000004fa_blk000004fb_sig0000157a,
      A1 => blk000004fa_blk000004fb_sig0000157b,
      A2 => blk000004fa_blk000004fb_sig0000157b,
      A3 => blk000004fa_blk000004fb_sig0000157b,
      CE => ce,
      CLK => clk,
      D => sig00000425,
      Q => blk000004fa_blk000004fb_sig00001583,
      Q15 => NLW_blk000004fa_blk000004fb_blk0000050c_Q15_UNCONNECTED
    );
  blk000004fa_blk000004fb_blk0000050b : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk000004fa_blk000004fb_sig00001582,
      Q => sig00000415
    );
  blk000004fa_blk000004fb_blk0000050a : SRLC16E
    generic map(
      INIT => X"0000"
    )
    port map (
      A0 => blk000004fa_blk000004fb_sig0000157a,
      A1 => blk000004fa_blk000004fb_sig0000157b,
      A2 => blk000004fa_blk000004fb_sig0000157b,
      A3 => blk000004fa_blk000004fb_sig0000157b,
      CE => ce,
      CLK => clk,
      D => sig00000423,
      Q => blk000004fa_blk000004fb_sig00001582,
      Q15 => NLW_blk000004fa_blk000004fb_blk0000050a_Q15_UNCONNECTED
    );
  blk000004fa_blk000004fb_blk00000509 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk000004fa_blk000004fb_sig00001581,
      Q => sig00000414
    );
  blk000004fa_blk000004fb_blk00000508 : SRLC16E
    generic map(
      INIT => X"0000"
    )
    port map (
      A0 => blk000004fa_blk000004fb_sig0000157a,
      A1 => blk000004fa_blk000004fb_sig0000157b,
      A2 => blk000004fa_blk000004fb_sig0000157b,
      A3 => blk000004fa_blk000004fb_sig0000157b,
      CE => ce,
      CLK => clk,
      D => sig00000422,
      Q => blk000004fa_blk000004fb_sig00001581,
      Q15 => NLW_blk000004fa_blk000004fb_blk00000508_Q15_UNCONNECTED
    );
  blk000004fa_blk000004fb_blk00000507 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk000004fa_blk000004fb_sig00001580,
      Q => sig00000416
    );
  blk000004fa_blk000004fb_blk00000506 : SRLC16E
    generic map(
      INIT => X"0000"
    )
    port map (
      A0 => blk000004fa_blk000004fb_sig0000157a,
      A1 => blk000004fa_blk000004fb_sig0000157b,
      A2 => blk000004fa_blk000004fb_sig0000157b,
      A3 => blk000004fa_blk000004fb_sig0000157b,
      CE => ce,
      CLK => clk,
      D => sig00000424,
      Q => blk000004fa_blk000004fb_sig00001580,
      Q15 => NLW_blk000004fa_blk000004fb_blk00000506_Q15_UNCONNECTED
    );
  blk000004fa_blk000004fb_blk00000505 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk000004fa_blk000004fb_sig0000157f,
      Q => sig00000413
    );
  blk000004fa_blk000004fb_blk00000504 : SRLC16E
    generic map(
      INIT => X"0000"
    )
    port map (
      A0 => blk000004fa_blk000004fb_sig0000157a,
      A1 => blk000004fa_blk000004fb_sig0000157b,
      A2 => blk000004fa_blk000004fb_sig0000157b,
      A3 => blk000004fa_blk000004fb_sig0000157b,
      CE => ce,
      CLK => clk,
      D => sig00000421,
      Q => blk000004fa_blk000004fb_sig0000157f,
      Q15 => NLW_blk000004fa_blk000004fb_blk00000504_Q15_UNCONNECTED
    );
  blk000004fa_blk000004fb_blk00000503 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk000004fa_blk000004fb_sig0000157e,
      Q => sig00000412
    );
  blk000004fa_blk000004fb_blk00000502 : SRLC16E
    generic map(
      INIT => X"0000"
    )
    port map (
      A0 => blk000004fa_blk000004fb_sig0000157a,
      A1 => blk000004fa_blk000004fb_sig0000157b,
      A2 => blk000004fa_blk000004fb_sig0000157b,
      A3 => blk000004fa_blk000004fb_sig0000157b,
      CE => ce,
      CLK => clk,
      D => sig00000420,
      Q => blk000004fa_blk000004fb_sig0000157e,
      Q15 => NLW_blk000004fa_blk000004fb_blk00000502_Q15_UNCONNECTED
    );
  blk000004fa_blk000004fb_blk00000501 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk000004fa_blk000004fb_sig0000157d,
      Q => sig00000411
    );
  blk000004fa_blk000004fb_blk00000500 : SRLC16E
    generic map(
      INIT => X"0000"
    )
    port map (
      A0 => blk000004fa_blk000004fb_sig0000157a,
      A1 => blk000004fa_blk000004fb_sig0000157b,
      A2 => blk000004fa_blk000004fb_sig0000157b,
      A3 => blk000004fa_blk000004fb_sig0000157b,
      CE => ce,
      CLK => clk,
      D => sig0000041f,
      Q => blk000004fa_blk000004fb_sig0000157d,
      Q15 => NLW_blk000004fa_blk000004fb_blk00000500_Q15_UNCONNECTED
    );
  blk000004fa_blk000004fb_blk000004ff : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk000004fa_blk000004fb_sig0000157c,
      Q => sig00000410
    );
  blk000004fa_blk000004fb_blk000004fe : SRLC16E
    generic map(
      INIT => X"0000"
    )
    port map (
      A0 => blk000004fa_blk000004fb_sig0000157a,
      A1 => blk000004fa_blk000004fb_sig0000157b,
      A2 => blk000004fa_blk000004fb_sig0000157b,
      A3 => blk000004fa_blk000004fb_sig0000157b,
      CE => ce,
      CLK => clk,
      D => sig0000041e,
      Q => blk000004fa_blk000004fb_sig0000157c,
      Q15 => NLW_blk000004fa_blk000004fb_blk000004fe_Q15_UNCONNECTED
    );
  blk000004fa_blk000004fb_blk000004fd : VCC
    port map (
      P => blk000004fa_blk000004fb_sig0000157b
    );
  blk000004fa_blk000004fb_blk000004fc : GND
    port map (
      G => blk000004fa_blk000004fb_sig0000157a
    );
  blk0000051a_blk0000051b_blk00000539 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk0000051a_blk0000051b_sig000015d6,
      Q => sig0000024d
    );
  blk0000051a_blk0000051b_blk00000538 : SRLC16E
    generic map(
      INIT => X"0000"
    )
    port map (
      A0 => blk0000051a_blk0000051b_sig000015c7,
      A1 => blk0000051a_blk0000051b_sig000015c8,
      A2 => blk0000051a_blk0000051b_sig000015c8,
      A3 => blk0000051a_blk0000051b_sig000015c8,
      CE => ce,
      CLK => clk,
      D => sig0000040e,
      Q => blk0000051a_blk0000051b_sig000015d6,
      Q15 => NLW_blk0000051a_blk0000051b_blk00000538_Q15_UNCONNECTED
    );
  blk0000051a_blk0000051b_blk00000537 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk0000051a_blk0000051b_sig000015d5,
      Q => sig0000024c
    );
  blk0000051a_blk0000051b_blk00000536 : SRLC16E
    generic map(
      INIT => X"0000"
    )
    port map (
      A0 => blk0000051a_blk0000051b_sig000015c7,
      A1 => blk0000051a_blk0000051b_sig000015c8,
      A2 => blk0000051a_blk0000051b_sig000015c8,
      A3 => blk0000051a_blk0000051b_sig000015c8,
      CE => ce,
      CLK => clk,
      D => sig0000040d,
      Q => blk0000051a_blk0000051b_sig000015d5,
      Q15 => NLW_blk0000051a_blk0000051b_blk00000536_Q15_UNCONNECTED
    );
  blk0000051a_blk0000051b_blk00000535 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk0000051a_blk0000051b_sig000015d4,
      Q => sig0000024e
    );
  blk0000051a_blk0000051b_blk00000534 : SRLC16E
    generic map(
      INIT => X"0000"
    )
    port map (
      A0 => blk0000051a_blk0000051b_sig000015c7,
      A1 => blk0000051a_blk0000051b_sig000015c8,
      A2 => blk0000051a_blk0000051b_sig000015c8,
      A3 => blk0000051a_blk0000051b_sig000015c8,
      CE => ce,
      CLK => clk,
      D => sig0000040f,
      Q => blk0000051a_blk0000051b_sig000015d4,
      Q15 => NLW_blk0000051a_blk0000051b_blk00000534_Q15_UNCONNECTED
    );
  blk0000051a_blk0000051b_blk00000533 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk0000051a_blk0000051b_sig000015d3,
      Q => sig0000024b
    );
  blk0000051a_blk0000051b_blk00000532 : SRLC16E
    generic map(
      INIT => X"0000"
    )
    port map (
      A0 => blk0000051a_blk0000051b_sig000015c7,
      A1 => blk0000051a_blk0000051b_sig000015c8,
      A2 => blk0000051a_blk0000051b_sig000015c8,
      A3 => blk0000051a_blk0000051b_sig000015c8,
      CE => ce,
      CLK => clk,
      D => sig0000040c,
      Q => blk0000051a_blk0000051b_sig000015d3,
      Q15 => NLW_blk0000051a_blk0000051b_blk00000532_Q15_UNCONNECTED
    );
  blk0000051a_blk0000051b_blk00000531 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk0000051a_blk0000051b_sig000015d2,
      Q => sig0000024a
    );
  blk0000051a_blk0000051b_blk00000530 : SRLC16E
    generic map(
      INIT => X"0000"
    )
    port map (
      A0 => blk0000051a_blk0000051b_sig000015c7,
      A1 => blk0000051a_blk0000051b_sig000015c8,
      A2 => blk0000051a_blk0000051b_sig000015c8,
      A3 => blk0000051a_blk0000051b_sig000015c8,
      CE => ce,
      CLK => clk,
      D => sig0000040b,
      Q => blk0000051a_blk0000051b_sig000015d2,
      Q15 => NLW_blk0000051a_blk0000051b_blk00000530_Q15_UNCONNECTED
    );
  blk0000051a_blk0000051b_blk0000052f : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk0000051a_blk0000051b_sig000015d1,
      Q => sig00000249
    );
  blk0000051a_blk0000051b_blk0000052e : SRLC16E
    generic map(
      INIT => X"0000"
    )
    port map (
      A0 => blk0000051a_blk0000051b_sig000015c7,
      A1 => blk0000051a_blk0000051b_sig000015c8,
      A2 => blk0000051a_blk0000051b_sig000015c8,
      A3 => blk0000051a_blk0000051b_sig000015c8,
      CE => ce,
      CLK => clk,
      D => sig0000040a,
      Q => blk0000051a_blk0000051b_sig000015d1,
      Q15 => NLW_blk0000051a_blk0000051b_blk0000052e_Q15_UNCONNECTED
    );
  blk0000051a_blk0000051b_blk0000052d : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk0000051a_blk0000051b_sig000015d0,
      Q => sig00000248
    );
  blk0000051a_blk0000051b_blk0000052c : SRLC16E
    generic map(
      INIT => X"0000"
    )
    port map (
      A0 => blk0000051a_blk0000051b_sig000015c7,
      A1 => blk0000051a_blk0000051b_sig000015c8,
      A2 => blk0000051a_blk0000051b_sig000015c8,
      A3 => blk0000051a_blk0000051b_sig000015c8,
      CE => ce,
      CLK => clk,
      D => sig00000409,
      Q => blk0000051a_blk0000051b_sig000015d0,
      Q15 => NLW_blk0000051a_blk0000051b_blk0000052c_Q15_UNCONNECTED
    );
  blk0000051a_blk0000051b_blk0000052b : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk0000051a_blk0000051b_sig000015cf,
      Q => sig00000246
    );
  blk0000051a_blk0000051b_blk0000052a : SRLC16E
    generic map(
      INIT => X"0000"
    )
    port map (
      A0 => blk0000051a_blk0000051b_sig000015c7,
      A1 => blk0000051a_blk0000051b_sig000015c8,
      A2 => blk0000051a_blk0000051b_sig000015c8,
      A3 => blk0000051a_blk0000051b_sig000015c8,
      CE => ce,
      CLK => clk,
      D => sig00000407,
      Q => blk0000051a_blk0000051b_sig000015cf,
      Q15 => NLW_blk0000051a_blk0000051b_blk0000052a_Q15_UNCONNECTED
    );
  blk0000051a_blk0000051b_blk00000529 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk0000051a_blk0000051b_sig000015ce,
      Q => sig00000245
    );
  blk0000051a_blk0000051b_blk00000528 : SRLC16E
    generic map(
      INIT => X"0000"
    )
    port map (
      A0 => blk0000051a_blk0000051b_sig000015c7,
      A1 => blk0000051a_blk0000051b_sig000015c8,
      A2 => blk0000051a_blk0000051b_sig000015c8,
      A3 => blk0000051a_blk0000051b_sig000015c8,
      CE => ce,
      CLK => clk,
      D => sig00000406,
      Q => blk0000051a_blk0000051b_sig000015ce,
      Q15 => NLW_blk0000051a_blk0000051b_blk00000528_Q15_UNCONNECTED
    );
  blk0000051a_blk0000051b_blk00000527 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk0000051a_blk0000051b_sig000015cd,
      Q => sig00000247
    );
  blk0000051a_blk0000051b_blk00000526 : SRLC16E
    generic map(
      INIT => X"0000"
    )
    port map (
      A0 => blk0000051a_blk0000051b_sig000015c7,
      A1 => blk0000051a_blk0000051b_sig000015c8,
      A2 => blk0000051a_blk0000051b_sig000015c8,
      A3 => blk0000051a_blk0000051b_sig000015c8,
      CE => ce,
      CLK => clk,
      D => sig00000408,
      Q => blk0000051a_blk0000051b_sig000015cd,
      Q15 => NLW_blk0000051a_blk0000051b_blk00000526_Q15_UNCONNECTED
    );
  blk0000051a_blk0000051b_blk00000525 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk0000051a_blk0000051b_sig000015cc,
      Q => sig00000244
    );
  blk0000051a_blk0000051b_blk00000524 : SRLC16E
    generic map(
      INIT => X"0000"
    )
    port map (
      A0 => blk0000051a_blk0000051b_sig000015c7,
      A1 => blk0000051a_blk0000051b_sig000015c8,
      A2 => blk0000051a_blk0000051b_sig000015c8,
      A3 => blk0000051a_blk0000051b_sig000015c8,
      CE => ce,
      CLK => clk,
      D => sig00000405,
      Q => blk0000051a_blk0000051b_sig000015cc,
      Q15 => NLW_blk0000051a_blk0000051b_blk00000524_Q15_UNCONNECTED
    );
  blk0000051a_blk0000051b_blk00000523 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk0000051a_blk0000051b_sig000015cb,
      Q => sig00000243
    );
  blk0000051a_blk0000051b_blk00000522 : SRLC16E
    generic map(
      INIT => X"0000"
    )
    port map (
      A0 => blk0000051a_blk0000051b_sig000015c7,
      A1 => blk0000051a_blk0000051b_sig000015c8,
      A2 => blk0000051a_blk0000051b_sig000015c8,
      A3 => blk0000051a_blk0000051b_sig000015c8,
      CE => ce,
      CLK => clk,
      D => sig00000404,
      Q => blk0000051a_blk0000051b_sig000015cb,
      Q15 => NLW_blk0000051a_blk0000051b_blk00000522_Q15_UNCONNECTED
    );
  blk0000051a_blk0000051b_blk00000521 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk0000051a_blk0000051b_sig000015ca,
      Q => sig00000242
    );
  blk0000051a_blk0000051b_blk00000520 : SRLC16E
    generic map(
      INIT => X"0000"
    )
    port map (
      A0 => blk0000051a_blk0000051b_sig000015c7,
      A1 => blk0000051a_blk0000051b_sig000015c8,
      A2 => blk0000051a_blk0000051b_sig000015c8,
      A3 => blk0000051a_blk0000051b_sig000015c8,
      CE => ce,
      CLK => clk,
      D => sig00000403,
      Q => blk0000051a_blk0000051b_sig000015ca,
      Q15 => NLW_blk0000051a_blk0000051b_blk00000520_Q15_UNCONNECTED
    );
  blk0000051a_blk0000051b_blk0000051f : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk0000051a_blk0000051b_sig000015c9,
      Q => sig00000241
    );
  blk0000051a_blk0000051b_blk0000051e : SRLC16E
    generic map(
      INIT => X"0000"
    )
    port map (
      A0 => blk0000051a_blk0000051b_sig000015c7,
      A1 => blk0000051a_blk0000051b_sig000015c8,
      A2 => blk0000051a_blk0000051b_sig000015c8,
      A3 => blk0000051a_blk0000051b_sig000015c8,
      CE => ce,
      CLK => clk,
      D => sig00000402,
      Q => blk0000051a_blk0000051b_sig000015c9,
      Q15 => NLW_blk0000051a_blk0000051b_blk0000051e_Q15_UNCONNECTED
    );
  blk0000051a_blk0000051b_blk0000051d : VCC
    port map (
      P => blk0000051a_blk0000051b_sig000015c8
    );
  blk0000051a_blk0000051b_blk0000051c : GND
    port map (
      G => blk0000051a_blk0000051b_sig000015c7
    );
  blk0000053a_blk00000572 : LUT2
    generic map(
      INIT => X"6"
    )
    port map (
      I0 => sig0000046d,
      I1 => sig00000443,
      O => blk0000053a_sig00001615
    );
  blk0000053a_blk00000571 : LUT2
    generic map(
      INIT => X"6"
    )
    port map (
      I0 => sig0000046c,
      I1 => sig00000442,
      O => blk0000053a_sig00001616
    );
  blk0000053a_blk00000570 : LUT2
    generic map(
      INIT => X"6"
    )
    port map (
      I0 => sig0000046b,
      I1 => sig00000441,
      O => blk0000053a_sig00001617
    );
  blk0000053a_blk0000056f : LUT2
    generic map(
      INIT => X"6"
    )
    port map (
      I0 => sig0000046a,
      I1 => sig00000440,
      O => blk0000053a_sig00001618
    );
  blk0000053a_blk0000056e : LUT2
    generic map(
      INIT => X"6"
    )
    port map (
      I0 => sig00000469,
      I1 => sig0000043f,
      O => blk0000053a_sig00001619
    );
  blk0000053a_blk0000056d : LUT2
    generic map(
      INIT => X"6"
    )
    port map (
      I0 => sig00000468,
      I1 => sig0000043e,
      O => blk0000053a_sig0000161a
    );
  blk0000053a_blk0000056c : LUT2
    generic map(
      INIT => X"6"
    )
    port map (
      I0 => sig00000467,
      I1 => sig0000043d,
      O => blk0000053a_sig0000161b
    );
  blk0000053a_blk0000056b : LUT2
    generic map(
      INIT => X"6"
    )
    port map (
      I0 => sig00000466,
      I1 => sig0000043c,
      O => blk0000053a_sig0000161c
    );
  blk0000053a_blk0000056a : LUT2
    generic map(
      INIT => X"6"
    )
    port map (
      I0 => sig00000465,
      I1 => sig0000043b,
      O => blk0000053a_sig0000161d
    );
  blk0000053a_blk00000569 : LUT2
    generic map(
      INIT => X"6"
    )
    port map (
      I0 => sig00000471,
      I1 => sig00000447,
      O => blk0000053a_sig0000161e
    );
  blk0000053a_blk00000568 : LUT2
    generic map(
      INIT => X"6"
    )
    port map (
      I0 => sig00000470,
      I1 => sig00000446,
      O => blk0000053a_sig00001612
    );
  blk0000053a_blk00000567 : LUT2
    generic map(
      INIT => X"6"
    )
    port map (
      I0 => sig0000046f,
      I1 => sig00000445,
      O => blk0000053a_sig00001613
    );
  blk0000053a_blk00000566 : LUT2
    generic map(
      INIT => X"6"
    )
    port map (
      I0 => sig0000046e,
      I1 => sig00000444,
      O => blk0000053a_sig00001614
    );
  blk0000053a_blk00000565 : LUT2
    generic map(
      INIT => X"6"
    )
    port map (
      I0 => sig00000464,
      I1 => sig0000043a,
      O => blk0000053a_sig0000161f
    );
  blk0000053a_blk00000564 : MUXCY
    port map (
      CI => blk0000053a_sig00001603,
      DI => sig00000464,
      S => blk0000053a_sig0000161f,
      O => blk0000053a_sig0000162c
    );
  blk0000053a_blk00000563 : MUXCY
    port map (
      CI => blk0000053a_sig0000162c,
      DI => sig00000465,
      S => blk0000053a_sig0000161d,
      O => blk0000053a_sig0000162b
    );
  blk0000053a_blk00000562 : MUXCY
    port map (
      CI => blk0000053a_sig0000162b,
      DI => sig00000466,
      S => blk0000053a_sig0000161c,
      O => blk0000053a_sig0000162a
    );
  blk0000053a_blk00000561 : MUXCY
    port map (
      CI => blk0000053a_sig0000162a,
      DI => sig00000467,
      S => blk0000053a_sig0000161b,
      O => blk0000053a_sig00001629
    );
  blk0000053a_blk00000560 : MUXCY
    port map (
      CI => blk0000053a_sig00001629,
      DI => sig00000468,
      S => blk0000053a_sig0000161a,
      O => blk0000053a_sig00001628
    );
  blk0000053a_blk0000055f : MUXCY
    port map (
      CI => blk0000053a_sig00001628,
      DI => sig00000469,
      S => blk0000053a_sig00001619,
      O => blk0000053a_sig00001627
    );
  blk0000053a_blk0000055e : MUXCY
    port map (
      CI => blk0000053a_sig00001627,
      DI => sig0000046a,
      S => blk0000053a_sig00001618,
      O => blk0000053a_sig00001626
    );
  blk0000053a_blk0000055d : MUXCY
    port map (
      CI => blk0000053a_sig00001626,
      DI => sig0000046b,
      S => blk0000053a_sig00001617,
      O => blk0000053a_sig00001625
    );
  blk0000053a_blk0000055c : MUXCY
    port map (
      CI => blk0000053a_sig00001625,
      DI => sig0000046c,
      S => blk0000053a_sig00001616,
      O => blk0000053a_sig00001624
    );
  blk0000053a_blk0000055b : MUXCY
    port map (
      CI => blk0000053a_sig00001624,
      DI => sig0000046d,
      S => blk0000053a_sig00001615,
      O => blk0000053a_sig00001623
    );
  blk0000053a_blk0000055a : MUXCY
    port map (
      CI => blk0000053a_sig00001623,
      DI => sig0000046e,
      S => blk0000053a_sig00001614,
      O => blk0000053a_sig00001622
    );
  blk0000053a_blk00000559 : MUXCY
    port map (
      CI => blk0000053a_sig00001622,
      DI => sig0000046f,
      S => blk0000053a_sig00001613,
      O => blk0000053a_sig00001621
    );
  blk0000053a_blk00000558 : MUXCY
    port map (
      CI => blk0000053a_sig00001621,
      DI => sig00000470,
      S => blk0000053a_sig00001612,
      O => blk0000053a_sig00001620
    );
  blk0000053a_blk00000557 : XORCY
    port map (
      CI => blk0000053a_sig00001603,
      LI => blk0000053a_sig0000161f,
      O => blk0000053a_sig00001611
    );
  blk0000053a_blk00000556 : XORCY
    port map (
      CI => blk0000053a_sig0000162c,
      LI => blk0000053a_sig0000161d,
      O => blk0000053a_sig00001610
    );
  blk0000053a_blk00000555 : XORCY
    port map (
      CI => blk0000053a_sig0000162b,
      LI => blk0000053a_sig0000161c,
      O => blk0000053a_sig0000160f
    );
  blk0000053a_blk00000554 : XORCY
    port map (
      CI => blk0000053a_sig0000162a,
      LI => blk0000053a_sig0000161b,
      O => blk0000053a_sig0000160e
    );
  blk0000053a_blk00000553 : XORCY
    port map (
      CI => blk0000053a_sig00001629,
      LI => blk0000053a_sig0000161a,
      O => blk0000053a_sig0000160d
    );
  blk0000053a_blk00000552 : XORCY
    port map (
      CI => blk0000053a_sig00001628,
      LI => blk0000053a_sig00001619,
      O => blk0000053a_sig0000160c
    );
  blk0000053a_blk00000551 : XORCY
    port map (
      CI => blk0000053a_sig00001627,
      LI => blk0000053a_sig00001618,
      O => blk0000053a_sig0000160b
    );
  blk0000053a_blk00000550 : XORCY
    port map (
      CI => blk0000053a_sig00001626,
      LI => blk0000053a_sig00001617,
      O => blk0000053a_sig0000160a
    );
  blk0000053a_blk0000054f : XORCY
    port map (
      CI => blk0000053a_sig00001625,
      LI => blk0000053a_sig00001616,
      O => blk0000053a_sig00001609
    );
  blk0000053a_blk0000054e : XORCY
    port map (
      CI => blk0000053a_sig00001624,
      LI => blk0000053a_sig00001615,
      O => blk0000053a_sig00001608
    );
  blk0000053a_blk0000054d : XORCY
    port map (
      CI => blk0000053a_sig00001623,
      LI => blk0000053a_sig00001614,
      O => blk0000053a_sig00001607
    );
  blk0000053a_blk0000054c : XORCY
    port map (
      CI => blk0000053a_sig00001622,
      LI => blk0000053a_sig00001613,
      O => blk0000053a_sig00001606
    );
  blk0000053a_blk0000054b : XORCY
    port map (
      CI => blk0000053a_sig00001621,
      LI => blk0000053a_sig00001612,
      O => blk0000053a_sig00001605
    );
  blk0000053a_blk0000054a : XORCY
    port map (
      CI => blk0000053a_sig00001620,
      LI => blk0000053a_sig0000161e,
      O => blk0000053a_sig00001604
    );
  blk0000053a_blk00000549 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk0000053a_sig00001604,
      Q => sig00000439
    );
  blk0000053a_blk00000548 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk0000053a_sig00001605,
      Q => sig00000438
    );
  blk0000053a_blk00000547 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk0000053a_sig00001606,
      Q => sig00000437
    );
  blk0000053a_blk00000546 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk0000053a_sig00001607,
      Q => sig00000436
    );
  blk0000053a_blk00000545 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk0000053a_sig00001608,
      Q => sig00000435
    );
  blk0000053a_blk00000544 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk0000053a_sig00001609,
      Q => sig00000434
    );
  blk0000053a_blk00000543 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk0000053a_sig0000160a,
      Q => sig00000433
    );
  blk0000053a_blk00000542 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk0000053a_sig0000160b,
      Q => sig00000432
    );
  blk0000053a_blk00000541 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk0000053a_sig0000160c,
      Q => sig00000431
    );
  blk0000053a_blk00000540 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk0000053a_sig0000160d,
      Q => sig00000430
    );
  blk0000053a_blk0000053f : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk0000053a_sig0000160e,
      Q => sig0000042f
    );
  blk0000053a_blk0000053e : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk0000053a_sig0000160f,
      Q => sig0000042e
    );
  blk0000053a_blk0000053d : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk0000053a_sig00001610,
      Q => sig0000042d
    );
  blk0000053a_blk0000053c : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk0000053a_sig00001611,
      Q => sig0000042c
    );
  blk0000053a_blk0000053b : GND
    port map (
      G => blk0000053a_sig00001603
    );
  blk00000573_blk000005ab : LUT2
    generic map(
      INIT => X"9"
    )
    port map (
      I0 => sig0000046d,
      I1 => sig00000443,
      O => blk00000573_sig0000166a
    );
  blk00000573_blk000005aa : LUT2
    generic map(
      INIT => X"9"
    )
    port map (
      I0 => sig0000046c,
      I1 => sig00000442,
      O => blk00000573_sig0000166b
    );
  blk00000573_blk000005a9 : LUT2
    generic map(
      INIT => X"9"
    )
    port map (
      I0 => sig0000046b,
      I1 => sig00000441,
      O => blk00000573_sig0000166c
    );
  blk00000573_blk000005a8 : LUT2
    generic map(
      INIT => X"9"
    )
    port map (
      I0 => sig0000046a,
      I1 => sig00000440,
      O => blk00000573_sig0000166d
    );
  blk00000573_blk000005a7 : LUT2
    generic map(
      INIT => X"9"
    )
    port map (
      I0 => sig00000469,
      I1 => sig0000043f,
      O => blk00000573_sig0000166e
    );
  blk00000573_blk000005a6 : LUT2
    generic map(
      INIT => X"9"
    )
    port map (
      I0 => sig00000468,
      I1 => sig0000043e,
      O => blk00000573_sig0000166f
    );
  blk00000573_blk000005a5 : LUT2
    generic map(
      INIT => X"9"
    )
    port map (
      I0 => sig00000467,
      I1 => sig0000043d,
      O => blk00000573_sig00001670
    );
  blk00000573_blk000005a4 : LUT2
    generic map(
      INIT => X"9"
    )
    port map (
      I0 => sig00000466,
      I1 => sig0000043c,
      O => blk00000573_sig00001671
    );
  blk00000573_blk000005a3 : LUT2
    generic map(
      INIT => X"9"
    )
    port map (
      I0 => sig00000465,
      I1 => sig0000043b,
      O => blk00000573_sig00001672
    );
  blk00000573_blk000005a2 : LUT2
    generic map(
      INIT => X"9"
    )
    port map (
      I0 => sig00000471,
      I1 => sig00000447,
      O => blk00000573_sig00001673
    );
  blk00000573_blk000005a1 : LUT2
    generic map(
      INIT => X"9"
    )
    port map (
      I0 => sig00000470,
      I1 => sig00000446,
      O => blk00000573_sig00001667
    );
  blk00000573_blk000005a0 : LUT2
    generic map(
      INIT => X"9"
    )
    port map (
      I0 => sig0000046f,
      I1 => sig00000445,
      O => blk00000573_sig00001668
    );
  blk00000573_blk0000059f : LUT2
    generic map(
      INIT => X"9"
    )
    port map (
      I0 => sig0000046e,
      I1 => sig00000444,
      O => blk00000573_sig00001669
    );
  blk00000573_blk0000059e : LUT2
    generic map(
      INIT => X"9"
    )
    port map (
      I0 => sig00000464,
      I1 => sig0000043a,
      O => blk00000573_sig00001674
    );
  blk00000573_blk0000059d : MUXCY
    port map (
      CI => blk00000573_sig00001682,
      DI => sig00000464,
      S => blk00000573_sig00001674,
      O => blk00000573_sig00001681
    );
  blk00000573_blk0000059c : MUXCY
    port map (
      CI => blk00000573_sig00001681,
      DI => sig00000465,
      S => blk00000573_sig00001672,
      O => blk00000573_sig00001680
    );
  blk00000573_blk0000059b : MUXCY
    port map (
      CI => blk00000573_sig00001680,
      DI => sig00000466,
      S => blk00000573_sig00001671,
      O => blk00000573_sig0000167f
    );
  blk00000573_blk0000059a : MUXCY
    port map (
      CI => blk00000573_sig0000167f,
      DI => sig00000467,
      S => blk00000573_sig00001670,
      O => blk00000573_sig0000167e
    );
  blk00000573_blk00000599 : MUXCY
    port map (
      CI => blk00000573_sig0000167e,
      DI => sig00000468,
      S => blk00000573_sig0000166f,
      O => blk00000573_sig0000167d
    );
  blk00000573_blk00000598 : MUXCY
    port map (
      CI => blk00000573_sig0000167d,
      DI => sig00000469,
      S => blk00000573_sig0000166e,
      O => blk00000573_sig0000167c
    );
  blk00000573_blk00000597 : MUXCY
    port map (
      CI => blk00000573_sig0000167c,
      DI => sig0000046a,
      S => blk00000573_sig0000166d,
      O => blk00000573_sig0000167b
    );
  blk00000573_blk00000596 : MUXCY
    port map (
      CI => blk00000573_sig0000167b,
      DI => sig0000046b,
      S => blk00000573_sig0000166c,
      O => blk00000573_sig0000167a
    );
  blk00000573_blk00000595 : MUXCY
    port map (
      CI => blk00000573_sig0000167a,
      DI => sig0000046c,
      S => blk00000573_sig0000166b,
      O => blk00000573_sig00001679
    );
  blk00000573_blk00000594 : MUXCY
    port map (
      CI => blk00000573_sig00001679,
      DI => sig0000046d,
      S => blk00000573_sig0000166a,
      O => blk00000573_sig00001678
    );
  blk00000573_blk00000593 : MUXCY
    port map (
      CI => blk00000573_sig00001678,
      DI => sig0000046e,
      S => blk00000573_sig00001669,
      O => blk00000573_sig00001677
    );
  blk00000573_blk00000592 : MUXCY
    port map (
      CI => blk00000573_sig00001677,
      DI => sig0000046f,
      S => blk00000573_sig00001668,
      O => blk00000573_sig00001676
    );
  blk00000573_blk00000591 : MUXCY
    port map (
      CI => blk00000573_sig00001676,
      DI => sig00000470,
      S => blk00000573_sig00001667,
      O => blk00000573_sig00001675
    );
  blk00000573_blk00000590 : XORCY
    port map (
      CI => blk00000573_sig00001682,
      LI => blk00000573_sig00001674,
      O => blk00000573_sig00001666
    );
  blk00000573_blk0000058f : XORCY
    port map (
      CI => blk00000573_sig00001681,
      LI => blk00000573_sig00001672,
      O => blk00000573_sig00001665
    );
  blk00000573_blk0000058e : XORCY
    port map (
      CI => blk00000573_sig00001680,
      LI => blk00000573_sig00001671,
      O => blk00000573_sig00001664
    );
  blk00000573_blk0000058d : XORCY
    port map (
      CI => blk00000573_sig0000167f,
      LI => blk00000573_sig00001670,
      O => blk00000573_sig00001663
    );
  blk00000573_blk0000058c : XORCY
    port map (
      CI => blk00000573_sig0000167e,
      LI => blk00000573_sig0000166f,
      O => blk00000573_sig00001662
    );
  blk00000573_blk0000058b : XORCY
    port map (
      CI => blk00000573_sig0000167d,
      LI => blk00000573_sig0000166e,
      O => blk00000573_sig00001661
    );
  blk00000573_blk0000058a : XORCY
    port map (
      CI => blk00000573_sig0000167c,
      LI => blk00000573_sig0000166d,
      O => blk00000573_sig00001660
    );
  blk00000573_blk00000589 : XORCY
    port map (
      CI => blk00000573_sig0000167b,
      LI => blk00000573_sig0000166c,
      O => blk00000573_sig0000165f
    );
  blk00000573_blk00000588 : XORCY
    port map (
      CI => blk00000573_sig0000167a,
      LI => blk00000573_sig0000166b,
      O => blk00000573_sig0000165e
    );
  blk00000573_blk00000587 : XORCY
    port map (
      CI => blk00000573_sig00001679,
      LI => blk00000573_sig0000166a,
      O => blk00000573_sig0000165d
    );
  blk00000573_blk00000586 : XORCY
    port map (
      CI => blk00000573_sig00001678,
      LI => blk00000573_sig00001669,
      O => blk00000573_sig0000165c
    );
  blk00000573_blk00000585 : XORCY
    port map (
      CI => blk00000573_sig00001677,
      LI => blk00000573_sig00001668,
      O => blk00000573_sig0000165b
    );
  blk00000573_blk00000584 : XORCY
    port map (
      CI => blk00000573_sig00001676,
      LI => blk00000573_sig00001667,
      O => blk00000573_sig0000165a
    );
  blk00000573_blk00000583 : XORCY
    port map (
      CI => blk00000573_sig00001675,
      LI => blk00000573_sig00001673,
      O => blk00000573_sig00001659
    );
  blk00000573_blk00000582 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000573_sig00001659,
      Q => sig0000042b
    );
  blk00000573_blk00000581 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000573_sig0000165a,
      Q => sig0000042a
    );
  blk00000573_blk00000580 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000573_sig0000165b,
      Q => sig00000429
    );
  blk00000573_blk0000057f : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000573_sig0000165c,
      Q => sig00000428
    );
  blk00000573_blk0000057e : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000573_sig0000165d,
      Q => sig00000427
    );
  blk00000573_blk0000057d : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000573_sig0000165e,
      Q => sig00000426
    );
  blk00000573_blk0000057c : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000573_sig0000165f,
      Q => sig00000425
    );
  blk00000573_blk0000057b : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000573_sig00001660,
      Q => sig00000424
    );
  blk00000573_blk0000057a : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000573_sig00001661,
      Q => sig00000423
    );
  blk00000573_blk00000579 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000573_sig00001662,
      Q => sig00000422
    );
  blk00000573_blk00000578 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000573_sig00001663,
      Q => sig00000421
    );
  blk00000573_blk00000577 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000573_sig00001664,
      Q => sig00000420
    );
  blk00000573_blk00000576 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000573_sig00001665,
      Q => sig0000041f
    );
  blk00000573_blk00000575 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000573_sig00001666,
      Q => sig0000041e
    );
  blk00000573_blk00000574 : VCC
    port map (
      P => blk00000573_sig00001682
    );
  blk000005ac_blk000005ad_blk000005bb : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk000005ac_blk000005ad_sig000016a6,
      Q => sig0000022d
    );
  blk000005ac_blk000005ad_blk000005ba : SRLC32E
    generic map(
      INIT => X"00000000"
    )
    port map (
      CLK => clk,
      D => sig00000280,
      CE => ce,
      Q => blk000005ac_blk000005ad_sig000016a6,
      Q31 => NLW_blk000005ac_blk000005ad_blk000005ba_Q31_UNCONNECTED,
      A(4) => blk000005ac_blk000005ad_sig000016a0,
      A(3) => blk000005ac_blk000005ad_sig0000169f,
      A(2) => blk000005ac_blk000005ad_sig0000169f,
      A(1) => blk000005ac_blk000005ad_sig000016a0,
      A(0) => blk000005ac_blk000005ad_sig000016a0
    );
  blk000005ac_blk000005ad_blk000005b9 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk000005ac_blk000005ad_sig000016a5,
      Q => sig00000232
    );
  blk000005ac_blk000005ad_blk000005b8 : SRLC32E
    generic map(
      INIT => X"00000000"
    )
    port map (
      CLK => clk,
      D => sig0000027f,
      CE => ce,
      Q => blk000005ac_blk000005ad_sig000016a5,
      Q31 => NLW_blk000005ac_blk000005ad_blk000005b8_Q31_UNCONNECTED,
      A(4) => blk000005ac_blk000005ad_sig000016a0,
      A(3) => blk000005ac_blk000005ad_sig0000169f,
      A(2) => blk000005ac_blk000005ad_sig0000169f,
      A(1) => blk000005ac_blk000005ad_sig000016a0,
      A(0) => blk000005ac_blk000005ad_sig000016a0
    );
  blk000005ac_blk000005ad_blk000005b7 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk000005ac_blk000005ad_sig000016a4,
      Q => sig0000022e
    );
  blk000005ac_blk000005ad_blk000005b6 : SRLC32E
    generic map(
      INIT => X"00000000"
    )
    port map (
      CLK => clk,
      D => sig00000281,
      CE => ce,
      Q => blk000005ac_blk000005ad_sig000016a4,
      Q31 => NLW_blk000005ac_blk000005ad_blk000005b6_Q31_UNCONNECTED,
      A(4) => blk000005ac_blk000005ad_sig000016a0,
      A(3) => blk000005ac_blk000005ad_sig0000169f,
      A(2) => blk000005ac_blk000005ad_sig0000169f,
      A(1) => blk000005ac_blk000005ad_sig000016a0,
      A(0) => blk000005ac_blk000005ad_sig000016a0
    );
  blk000005ac_blk000005ad_blk000005b5 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk000005ac_blk000005ad_sig000016a3,
      Q => sig00000230
    );
  blk000005ac_blk000005ad_blk000005b4 : SRLC32E
    generic map(
      INIT => X"00000000"
    )
    port map (
      CLK => clk,
      D => sig0000027d,
      CE => ce,
      Q => blk000005ac_blk000005ad_sig000016a3,
      Q31 => NLW_blk000005ac_blk000005ad_blk000005b4_Q31_UNCONNECTED,
      A(4) => blk000005ac_blk000005ad_sig000016a0,
      A(3) => blk000005ac_blk000005ad_sig0000169f,
      A(2) => blk000005ac_blk000005ad_sig0000169f,
      A(1) => blk000005ac_blk000005ad_sig000016a0,
      A(0) => blk000005ac_blk000005ad_sig000016a0
    );
  blk000005ac_blk000005ad_blk000005b3 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk000005ac_blk000005ad_sig000016a2,
      Q => sig0000022f
    );
  blk000005ac_blk000005ad_blk000005b2 : SRLC32E
    generic map(
      INIT => X"00000000"
    )
    port map (
      CLK => clk,
      D => sig0000027c,
      CE => ce,
      Q => blk000005ac_blk000005ad_sig000016a2,
      Q31 => NLW_blk000005ac_blk000005ad_blk000005b2_Q31_UNCONNECTED,
      A(4) => blk000005ac_blk000005ad_sig000016a0,
      A(3) => blk000005ac_blk000005ad_sig0000169f,
      A(2) => blk000005ac_blk000005ad_sig0000169f,
      A(1) => blk000005ac_blk000005ad_sig000016a0,
      A(0) => blk000005ac_blk000005ad_sig000016a0
    );
  blk000005ac_blk000005ad_blk000005b1 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk000005ac_blk000005ad_sig000016a1,
      Q => sig00000231
    );
  blk000005ac_blk000005ad_blk000005b0 : SRLC32E
    generic map(
      INIT => X"00000000"
    )
    port map (
      CLK => clk,
      D => sig0000027e,
      CE => ce,
      Q => blk000005ac_blk000005ad_sig000016a1,
      Q31 => NLW_blk000005ac_blk000005ad_blk000005b0_Q31_UNCONNECTED,
      A(4) => blk000005ac_blk000005ad_sig000016a0,
      A(3) => blk000005ac_blk000005ad_sig0000169f,
      A(2) => blk000005ac_blk000005ad_sig0000169f,
      A(1) => blk000005ac_blk000005ad_sig000016a0,
      A(0) => blk000005ac_blk000005ad_sig000016a0
    );
  blk000005ac_blk000005ad_blk000005af : VCC
    port map (
      P => blk000005ac_blk000005ad_sig000016a0
    );
  blk000005ac_blk000005ad_blk000005ae : GND
    port map (
      G => blk000005ac_blk000005ad_sig0000169f
    );
  blk000005bc_blk000005bd_blk000005c1 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk000005bc_blk000005bd_sig000016b1,
      Q => sig0000022c
    );
  blk000005bc_blk000005bd_blk000005c0 : SRLC32E
    generic map(
      INIT => X"00000000"
    )
    port map (
      CLK => clk,
      D => sig000001eb,
      CE => ce,
      Q => blk000005bc_blk000005bd_sig000016b1,
      Q31 => NLW_blk000005bc_blk000005bd_blk000005c0_Q31_UNCONNECTED,
      A(4) => blk000005bc_blk000005bd_sig000016b0,
      A(3) => blk000005bc_blk000005bd_sig000016af,
      A(2) => blk000005bc_blk000005bd_sig000016af,
      A(1) => blk000005bc_blk000005bd_sig000016b0,
      A(0) => blk000005bc_blk000005bd_sig000016b0
    );
  blk000005bc_blk000005bd_blk000005bf : VCC
    port map (
      P => blk000005bc_blk000005bd_sig000016b0
    );
  blk000005bc_blk000005bd_blk000005be : GND
    port map (
      G => blk000005bc_blk000005bd_sig000016af
    );
  blk000005c2_blk000005c3_blk000005c6 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk000005c2_blk000005c3_sig000016c2,
      Q => sig00000497
    );
  blk000005c2_blk000005c3_blk000005c5 : SRLC16E
    generic map(
      INIT => X"0000"
    )
    port map (
      A0 => blk000005c2_blk000005c3_sig000016c1,
      A1 => blk000005c2_blk000005c3_sig000016c1,
      A2 => blk000005c2_blk000005c3_sig000016c1,
      A3 => blk000005c2_blk000005c3_sig000016c1,
      CE => ce,
      CLK => clk,
      D => sig00000498,
      Q => blk000005c2_blk000005c3_sig000016c2,
      Q15 => NLW_blk000005c2_blk000005c3_blk000005c5_Q15_UNCONNECTED
    );
  blk000005c2_blk000005c3_blk000005c4 : GND
    port map (
      G => blk000005c2_blk000005c3_sig000016c1
    );
  blk000005cd_blk000005e4 : LUT1
    generic map(
      INIT => X"2"
    )
    port map (
      I0 => sig0000022f,
      O => blk000005cd_sig000016e4
    );
  blk000005cd_blk000005e3 : LUT1
    generic map(
      INIT => X"2"
    )
    port map (
      I0 => sig00000232,
      O => blk000005cd_sig000016e3
    );
  blk000005cd_blk000005e2 : LUT2
    generic map(
      INIT => X"6"
    )
    port map (
      I0 => sig00000231,
      I1 => sig00000232,
      O => blk000005cd_sig000016db
    );
  blk000005cd_blk000005e1 : LUT2
    generic map(
      INIT => X"6"
    )
    port map (
      I0 => sig00000230,
      I1 => sig00000231,
      O => blk000005cd_sig000016dc
    );
  blk000005cd_blk000005e0 : LUT2
    generic map(
      INIT => X"6"
    )
    port map (
      I0 => sig0000022f,
      I1 => sig00000230,
      O => blk000005cd_sig000016dd
    );
  blk000005cd_blk000005df : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk000005cd_sig000016d5,
      Q => sig0000049e
    );
  blk000005cd_blk000005de : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk000005cd_sig000016da,
      Q => sig0000049f
    );
  blk000005cd_blk000005dd : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk000005cd_sig000016d9,
      Q => sig000004a0
    );
  blk000005cd_blk000005dc : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk000005cd_sig000016d8,
      Q => sig000004a1
    );
  blk000005cd_blk000005db : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk000005cd_sig000016d7,
      Q => sig000004a2
    );
  blk000005cd_blk000005da : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk000005cd_sig000016d6,
      Q => sig000004a3
    );
  blk000005cd_blk000005d9 : MUXCY
    port map (
      CI => blk000005cd_sig000016d4,
      DI => sig000008b6,
      S => blk000005cd_sig000016e4,
      O => blk000005cd_sig000016e2
    );
  blk000005cd_blk000005d8 : MUXCY
    port map (
      CI => blk000005cd_sig000016e2,
      DI => sig0000022f,
      S => blk000005cd_sig000016dd,
      O => blk000005cd_sig000016e1
    );
  blk000005cd_blk000005d7 : MUXCY
    port map (
      CI => blk000005cd_sig000016e1,
      DI => sig00000230,
      S => blk000005cd_sig000016dc,
      O => blk000005cd_sig000016e0
    );
  blk000005cd_blk000005d6 : MUXCY
    port map (
      CI => blk000005cd_sig000016e0,
      DI => sig00000231,
      S => blk000005cd_sig000016db,
      O => blk000005cd_sig000016df
    );
  blk000005cd_blk000005d5 : MUXCY
    port map (
      CI => blk000005cd_sig000016df,
      DI => sig00000232,
      S => blk000005cd_sig000016e3,
      O => blk000005cd_sig000016de
    );
  blk000005cd_blk000005d4 : XORCY
    port map (
      CI => blk000005cd_sig000016e2,
      LI => blk000005cd_sig000016dd,
      O => blk000005cd_sig000016da
    );
  blk000005cd_blk000005d3 : XORCY
    port map (
      CI => blk000005cd_sig000016e1,
      LI => blk000005cd_sig000016dc,
      O => blk000005cd_sig000016d9
    );
  blk000005cd_blk000005d2 : XORCY
    port map (
      CI => blk000005cd_sig000016e0,
      LI => blk000005cd_sig000016db,
      O => blk000005cd_sig000016d8
    );
  blk000005cd_blk000005d1 : XORCY
    port map (
      CI => blk000005cd_sig000016df,
      LI => blk000005cd_sig000016e3,
      O => blk000005cd_sig000016d7
    );
  blk000005cd_blk000005d0 : XORCY
    port map (
      CI => blk000005cd_sig000016de,
      LI => blk000005cd_sig000016d4,
      O => blk000005cd_sig000016d6
    );
  blk000005cd_blk000005cf : XORCY
    port map (
      CI => blk000005cd_sig000016d4,
      LI => blk000005cd_sig000016e4,
      O => blk000005cd_sig000016d5
    );
  blk000005cd_blk000005ce : GND
    port map (
      G => blk000005cd_sig000016d4
    );
  blk000005f1_blk00000654 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk000005f1_sig0000174f,
      Q => sig00000496
    );
  blk000005f1_blk00000653 : SRLC16E
    generic map(
      INIT => X"0000"
    )
    port map (
      A0 => blk000005f1_sig0000174e,
      A1 => blk000005f1_sig0000174e,
      A2 => blk000005f1_sig0000174e,
      A3 => blk000005f1_sig0000174e,
      CE => ce,
      CLK => clk,
      D => sig00000494,
      Q => blk000005f1_sig0000174f,
      Q15 => NLW_blk000005f1_blk00000653_Q15_UNCONNECTED
    );
  blk000005f1_blk00000652 : GND
    port map (
      G => blk000005f1_sig0000174e
    );
  blk000005f1_blk00000651 : LUT4
    generic map(
      INIT => X"AE28"
    )
    port map (
      I0 => sig0000049a,
      I1 => sig0000049c,
      I2 => sig0000049b,
      I3 => sig00000499,
      O => blk000005f1_sig00001738
    );
  blk000005f1_blk00000650 : LUT4
    generic map(
      INIT => X"A628"
    )
    port map (
      I0 => sig0000049c,
      I1 => sig0000049b,
      I2 => sig0000049a,
      I3 => sig00000499,
      O => blk000005f1_sig00001739
    );
  blk000005f1_blk0000064f : LUT4
    generic map(
      INIT => X"2B82"
    )
    port map (
      I0 => sig0000049c,
      I1 => sig0000049b,
      I2 => sig0000049a,
      I3 => sig00000499,
      O => blk000005f1_sig0000173a
    );
  blk000005f1_blk0000064e : LUT4
    generic map(
      INIT => X"86AA"
    )
    port map (
      I0 => sig0000049c,
      I1 => sig0000049b,
      I2 => sig00000499,
      I3 => sig0000049a,
      O => blk000005f1_sig0000173c
    );
  blk000005f1_blk0000064d : LUT4
    generic map(
      INIT => X"9A38"
    )
    port map (
      I0 => sig0000049b,
      I1 => sig0000049c,
      I2 => sig00000499,
      I3 => sig0000049a,
      O => blk000005f1_sig0000173d
    );
  blk000005f1_blk0000064c : LUT4
    generic map(
      INIT => X"EA44"
    )
    port map (
      I0 => sig0000049c,
      I1 => sig0000049a,
      I2 => sig0000049b,
      I3 => sig00000499,
      O => blk000005f1_sig00001742
    );
  blk000005f1_blk0000064b : LUT4
    generic map(
      INIT => X"7528"
    )
    port map (
      I0 => sig0000049a,
      I1 => sig0000049c,
      I2 => sig0000049b,
      I3 => sig00000499,
      O => blk000005f1_sig00001743
    );
  blk000005f1_blk0000064a : LUT4
    generic map(
      INIT => X"D142"
    )
    port map (
      I0 => sig0000049c,
      I1 => sig0000049b,
      I2 => sig00000499,
      I3 => sig0000049a,
      O => blk000005f1_sig00001745
    );
  blk000005f1_blk00000649 : LUT4
    generic map(
      INIT => X"A394"
    )
    port map (
      I0 => sig0000049c,
      I1 => sig0000049b,
      I2 => sig00000499,
      I3 => sig0000049a,
      O => blk000005f1_sig00001748
    );
  blk000005f1_blk00000648 : LUT4
    generic map(
      INIT => X"D1B4"
    )
    port map (
      I0 => sig0000049b,
      I1 => sig0000049c,
      I2 => sig0000049a,
      I3 => sig00000499,
      O => blk000005f1_sig00001749
    );
  blk000005f1_blk00000647 : LUT4
    generic map(
      INIT => X"657E"
    )
    port map (
      I0 => sig0000049b,
      I1 => sig00000499,
      I2 => sig0000049c,
      I3 => sig0000049a,
      O => blk000005f1_sig0000174a
    );
  blk000005f1_blk00000646 : LUT4
    generic map(
      INIT => X"8BD2"
    )
    port map (
      I0 => sig0000049c,
      I1 => sig0000049b,
      I2 => sig00000499,
      I3 => sig0000049a,
      O => blk000005f1_sig0000173e
    );
  blk000005f1_blk00000645 : LUT4
    generic map(
      INIT => X"5616"
    )
    port map (
      I0 => sig0000049c,
      I1 => sig0000049b,
      I2 => sig00000499,
      I3 => sig0000049a,
      O => blk000005f1_sig00001747
    );
  blk000005f1_blk00000644 : LUT4
    generic map(
      INIT => X"0BB8"
    )
    port map (
      I0 => sig0000049c,
      I1 => sig0000049b,
      I2 => sig0000049a,
      I3 => sig00000499,
      O => blk000005f1_sig00001746
    );
  blk000005f1_blk00000643 : LUT4
    generic map(
      INIT => X"EC9E"
    )
    port map (
      I0 => sig0000049c,
      I1 => sig0000049b,
      I2 => sig0000049a,
      I3 => sig00000499,
      O => blk000005f1_sig0000173f
    );
  blk000005f1_blk00000642 : LUT4
    generic map(
      INIT => X"0001"
    )
    port map (
      I0 => sig0000049c,
      I1 => sig0000049b,
      I2 => sig0000049a,
      I3 => sig00000499,
      O => blk000005f1_sig0000174d
    );
  blk000005f1_blk00000641 : LUT4
    generic map(
      INIT => X"557E"
    )
    port map (
      I0 => sig0000049c,
      I1 => sig00000499,
      I2 => sig0000049a,
      I3 => sig0000049b,
      O => blk000005f1_sig0000174c
    );
  blk000005f1_blk00000640 : LUT4
    generic map(
      INIT => X"BBE8"
    )
    port map (
      I0 => sig0000049c,
      I1 => sig0000049a,
      I2 => sig00000499,
      I3 => sig0000049b,
      O => blk000005f1_sig00001740
    );
  blk000005f1_blk0000063f : LUT4
    generic map(
      INIT => X"77D4"
    )
    port map (
      I0 => sig0000049c,
      I1 => sig0000049a,
      I2 => sig00000499,
      I3 => sig0000049b,
      O => blk000005f1_sig0000174b
    );
  blk000005f1_blk0000063e : LUT4
    generic map(
      INIT => X"8A8E"
    )
    port map (
      I0 => sig0000049a,
      I1 => sig0000049b,
      I2 => sig0000049c,
      I3 => sig00000499,
      O => blk000005f1_sig0000173b
    );
  blk000005f1_blk0000063d : LUT4
    generic map(
      INIT => X"626A"
    )
    port map (
      I0 => sig00000499,
      I1 => sig0000049c,
      I2 => sig0000049a,
      I3 => sig0000049b,
      O => blk000005f1_sig00001737
    );
  blk000005f1_blk0000063c : LUT4
    generic map(
      INIT => X"5584"
    )
    port map (
      I0 => sig0000049c,
      I1 => sig00000499,
      I2 => sig0000049a,
      I3 => sig0000049b,
      O => blk000005f1_sig00001744
    );
  blk000005f1_blk0000063b : LUT3
    generic map(
      INIT => X"D8"
    )
    port map (
      I0 => blk000005f1_sig000016f9,
      I1 => blk000005f1_sig0000171e,
      I2 => blk000005f1_sig000016f8,
      O => blk000005f1_sig00001736
    );
  blk000005f1_blk0000063a : LUT3
    generic map(
      INIT => X"D8"
    )
    port map (
      I0 => blk000005f1_sig000016f9,
      I1 => blk000005f1_sig00001714,
      I2 => blk000005f1_sig000016ee,
      O => blk000005f1_sig0000172c
    );
  blk000005f1_blk00000639 : LUT2
    generic map(
      INIT => X"4"
    )
    port map (
      I0 => blk000005f1_sig000016f9,
      I1 => blk000005f1_sig000016ed,
      O => blk000005f1_sig0000172b
    );
  blk000005f1_blk00000638 : LUT3
    generic map(
      INIT => X"D8"
    )
    port map (
      I0 => blk000005f1_sig000016f9,
      I1 => blk000005f1_sig0000171d,
      I2 => blk000005f1_sig000016f7,
      O => blk000005f1_sig00001735
    );
  blk000005f1_blk00000637 : LUT3
    generic map(
      INIT => X"D8"
    )
    port map (
      I0 => blk000005f1_sig000016f9,
      I1 => blk000005f1_sig0000171c,
      I2 => blk000005f1_sig000016f6,
      O => blk000005f1_sig00001734
    );
  blk000005f1_blk00000636 : LUT3
    generic map(
      INIT => X"D8"
    )
    port map (
      I0 => blk000005f1_sig000016f9,
      I1 => blk000005f1_sig0000171b,
      I2 => blk000005f1_sig000016f5,
      O => blk000005f1_sig00001733
    );
  blk000005f1_blk00000635 : LUT3
    generic map(
      INIT => X"D8"
    )
    port map (
      I0 => blk000005f1_sig000016f9,
      I1 => blk000005f1_sig0000171a,
      I2 => blk000005f1_sig000016f4,
      O => blk000005f1_sig00001732
    );
  blk000005f1_blk00000634 : LUT3
    generic map(
      INIT => X"D8"
    )
    port map (
      I0 => blk000005f1_sig000016f9,
      I1 => blk000005f1_sig00001719,
      I2 => blk000005f1_sig000016f3,
      O => blk000005f1_sig00001731
    );
  blk000005f1_blk00000633 : LUT3
    generic map(
      INIT => X"D8"
    )
    port map (
      I0 => blk000005f1_sig000016f9,
      I1 => blk000005f1_sig00001718,
      I2 => blk000005f1_sig000016f2,
      O => blk000005f1_sig00001730
    );
  blk000005f1_blk00000632 : LUT3
    generic map(
      INIT => X"D8"
    )
    port map (
      I0 => blk000005f1_sig000016f9,
      I1 => blk000005f1_sig00001717,
      I2 => blk000005f1_sig000016f1,
      O => blk000005f1_sig0000172f
    );
  blk000005f1_blk00000631 : LUT3
    generic map(
      INIT => X"D8"
    )
    port map (
      I0 => blk000005f1_sig000016f9,
      I1 => blk000005f1_sig00001716,
      I2 => blk000005f1_sig000016f0,
      O => blk000005f1_sig0000172e
    );
  blk000005f1_blk00000630 : LUT3
    generic map(
      INIT => X"D8"
    )
    port map (
      I0 => blk000005f1_sig000016f9,
      I1 => blk000005f1_sig00001715,
      I2 => blk000005f1_sig000016ef,
      O => blk000005f1_sig0000172d
    );
  blk000005f1_blk0000062f : LUT3
    generic map(
      INIT => X"D8"
    )
    port map (
      I0 => blk000005f1_sig000016f9,
      I1 => blk000005f1_sig000016f8,
      I2 => blk000005f1_sig0000171e,
      O => blk000005f1_sig0000172a
    );
  blk000005f1_blk0000062e : LUT3
    generic map(
      INIT => X"D8"
    )
    port map (
      I0 => blk000005f1_sig000016f9,
      I1 => blk000005f1_sig000016ee,
      I2 => blk000005f1_sig00001714,
      O => blk000005f1_sig00001720
    );
  blk000005f1_blk0000062d : LUT2
    generic map(
      INIT => X"8"
    )
    port map (
      I0 => blk000005f1_sig000016f9,
      I1 => blk000005f1_sig000016ed,
      O => blk000005f1_sig0000171f
    );
  blk000005f1_blk0000062c : LUT3
    generic map(
      INIT => X"D8"
    )
    port map (
      I0 => blk000005f1_sig000016f9,
      I1 => blk000005f1_sig000016f7,
      I2 => blk000005f1_sig0000171d,
      O => blk000005f1_sig00001729
    );
  blk000005f1_blk0000062b : LUT3
    generic map(
      INIT => X"D8"
    )
    port map (
      I0 => blk000005f1_sig000016f9,
      I1 => blk000005f1_sig000016f6,
      I2 => blk000005f1_sig0000171c,
      O => blk000005f1_sig00001728
    );
  blk000005f1_blk0000062a : LUT3
    generic map(
      INIT => X"D8"
    )
    port map (
      I0 => blk000005f1_sig000016f9,
      I1 => blk000005f1_sig000016f5,
      I2 => blk000005f1_sig0000171b,
      O => blk000005f1_sig00001727
    );
  blk000005f1_blk00000629 : LUT3
    generic map(
      INIT => X"D8"
    )
    port map (
      I0 => blk000005f1_sig000016f9,
      I1 => blk000005f1_sig000016f4,
      I2 => blk000005f1_sig0000171a,
      O => blk000005f1_sig00001726
    );
  blk000005f1_blk00000628 : LUT3
    generic map(
      INIT => X"D8"
    )
    port map (
      I0 => blk000005f1_sig000016f9,
      I1 => blk000005f1_sig000016f3,
      I2 => blk000005f1_sig00001719,
      O => blk000005f1_sig00001725
    );
  blk000005f1_blk00000627 : LUT3
    generic map(
      INIT => X"D8"
    )
    port map (
      I0 => blk000005f1_sig000016f9,
      I1 => blk000005f1_sig000016f2,
      I2 => blk000005f1_sig00001718,
      O => blk000005f1_sig00001724
    );
  blk000005f1_blk00000626 : LUT3
    generic map(
      INIT => X"D8"
    )
    port map (
      I0 => blk000005f1_sig000016f9,
      I1 => blk000005f1_sig000016f1,
      I2 => blk000005f1_sig00001717,
      O => blk000005f1_sig00001723
    );
  blk000005f1_blk00000625 : LUT3
    generic map(
      INIT => X"D8"
    )
    port map (
      I0 => blk000005f1_sig000016f9,
      I1 => blk000005f1_sig000016f0,
      I2 => blk000005f1_sig00001716,
      O => blk000005f1_sig00001722
    );
  blk000005f1_blk00000624 : LUT3
    generic map(
      INIT => X"D8"
    )
    port map (
      I0 => blk000005f1_sig000016f9,
      I1 => blk000005f1_sig000016ef,
      I2 => blk000005f1_sig00001715,
      O => blk000005f1_sig00001721
    );
  blk000005f1_blk00000623 : LUT3
    generic map(
      INIT => X"F8"
    )
    port map (
      I0 => sig0000049a,
      I1 => sig0000049b,
      I2 => sig0000049c,
      O => blk000005f1_sig00001741
    );
  blk000005f1_blk00000622 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk000005f1_sig0000172b,
      Q => sig0000022b
    );
  blk000005f1_blk00000621 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk000005f1_sig0000172c,
      Q => sig0000022a
    );
  blk000005f1_blk00000620 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk000005f1_sig0000172d,
      Q => sig00000229
    );
  blk000005f1_blk0000061f : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk000005f1_sig0000172e,
      Q => sig00000228
    );
  blk000005f1_blk0000061e : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk000005f1_sig0000172f,
      Q => sig00000227
    );
  blk000005f1_blk0000061d : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk000005f1_sig00001730,
      Q => sig00000226
    );
  blk000005f1_blk0000061c : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk000005f1_sig00001731,
      Q => sig00000225
    );
  blk000005f1_blk0000061b : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk000005f1_sig00001732,
      Q => sig00000224
    );
  blk000005f1_blk0000061a : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk000005f1_sig00001733,
      Q => sig00000223
    );
  blk000005f1_blk00000619 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk000005f1_sig00001734,
      Q => sig00000222
    );
  blk000005f1_blk00000618 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk000005f1_sig00001735,
      Q => sig00000221
    );
  blk000005f1_blk00000617 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk000005f1_sig00001736,
      Q => sig00000220
    );
  blk000005f1_blk00000616 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk000005f1_sig0000171f,
      Q => sig0000021f
    );
  blk000005f1_blk00000615 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk000005f1_sig00001720,
      Q => sig0000021e
    );
  blk000005f1_blk00000614 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk000005f1_sig00001721,
      Q => sig0000021d
    );
  blk000005f1_blk00000613 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk000005f1_sig00001722,
      Q => sig0000021c
    );
  blk000005f1_blk00000612 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk000005f1_sig00001723,
      Q => sig0000021b
    );
  blk000005f1_blk00000611 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk000005f1_sig00001724,
      Q => sig0000021a
    );
  blk000005f1_blk00000610 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk000005f1_sig00001725,
      Q => sig00000219
    );
  blk000005f1_blk0000060f : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk000005f1_sig00001726,
      Q => sig00000218
    );
  blk000005f1_blk0000060e : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk000005f1_sig00001727,
      Q => sig00000217
    );
  blk000005f1_blk0000060d : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk000005f1_sig00001728,
      Q => sig00000216
    );
  blk000005f1_blk0000060c : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk000005f1_sig00001729,
      Q => sig00000215
    );
  blk000005f1_blk0000060b : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk000005f1_sig0000172a,
      Q => sig00000214
    );
  blk000005f1_blk0000060a : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk000005f1_sig00001741,
      Q => blk000005f1_sig00001714
    );
  blk000005f1_blk00000609 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk000005f1_sig00001740,
      Q => blk000005f1_sig00001715
    );
  blk000005f1_blk00000608 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk000005f1_sig0000173f,
      Q => blk000005f1_sig00001716
    );
  blk000005f1_blk00000607 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk000005f1_sig0000173e,
      Q => blk000005f1_sig00001717
    );
  blk000005f1_blk00000606 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk000005f1_sig0000173d,
      Q => blk000005f1_sig00001718
    );
  blk000005f1_blk00000605 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk000005f1_sig0000173c,
      Q => blk000005f1_sig00001719
    );
  blk000005f1_blk00000604 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk000005f1_sig0000173b,
      Q => blk000005f1_sig0000171a
    );
  blk000005f1_blk00000603 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk000005f1_sig0000173a,
      Q => blk000005f1_sig0000171b
    );
  blk000005f1_blk00000602 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk000005f1_sig00001739,
      Q => blk000005f1_sig0000171c
    );
  blk000005f1_blk00000601 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk000005f1_sig00001738,
      Q => blk000005f1_sig0000171d
    );
  blk000005f1_blk00000600 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk000005f1_sig00001737,
      Q => blk000005f1_sig0000171e
    );
  blk000005f1_blk000005ff : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk000005f1_sig000016f9,
      Q => sig00000495
    );
  blk000005f1_blk000005fe : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk000005f1_sig0000174d,
      Q => blk000005f1_sig000016ed
    );
  blk000005f1_blk000005fd : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk000005f1_sig0000174c,
      Q => blk000005f1_sig000016ee
    );
  blk000005f1_blk000005fc : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk000005f1_sig0000174b,
      Q => blk000005f1_sig000016ef
    );
  blk000005f1_blk000005fb : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk000005f1_sig0000174a,
      Q => blk000005f1_sig000016f0
    );
  blk000005f1_blk000005fa : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk000005f1_sig00001749,
      Q => blk000005f1_sig000016f1
    );
  blk000005f1_blk000005f9 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk000005f1_sig00001748,
      Q => blk000005f1_sig000016f2
    );
  blk000005f1_blk000005f8 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk000005f1_sig00001747,
      Q => blk000005f1_sig000016f3
    );
  blk000005f1_blk000005f7 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk000005f1_sig00001746,
      Q => blk000005f1_sig000016f4
    );
  blk000005f1_blk000005f6 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk000005f1_sig00001745,
      Q => blk000005f1_sig000016f5
    );
  blk000005f1_blk000005f5 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk000005f1_sig00001744,
      Q => blk000005f1_sig000016f6
    );
  blk000005f1_blk000005f4 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk000005f1_sig00001743,
      Q => blk000005f1_sig000016f7
    );
  blk000005f1_blk000005f3 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk000005f1_sig00001742,
      Q => blk000005f1_sig000016f8
    );
  blk000005f1_blk000005f2 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => sig0000049d,
      Q => blk000005f1_sig000016f9
    );
  blk0000091a_blk0000091b_blk0000091f : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk0000091a_blk0000091b_sig0000195f,
      Q => sig00000a36
    );
  blk0000091a_blk0000091b_blk0000091e : SRLC16E
    generic map(
      INIT => X"0000"
    )
    port map (
      A0 => blk0000091a_blk0000091b_sig0000195d,
      A1 => blk0000091a_blk0000091b_sig0000195e,
      A2 => blk0000091a_blk0000091b_sig0000195e,
      A3 => blk0000091a_blk0000091b_sig0000195e,
      CE => ce,
      CLK => clk,
      D => sig000009f9,
      Q => blk0000091a_blk0000091b_sig0000195f,
      Q15 => NLW_blk0000091a_blk0000091b_blk0000091e_Q15_UNCONNECTED
    );
  blk0000091a_blk0000091b_blk0000091d : VCC
    port map (
      P => blk0000091a_blk0000091b_sig0000195e
    );
  blk0000091a_blk0000091b_blk0000091c : GND
    port map (
      G => blk0000091a_blk0000091b_sig0000195d
    );
  blk0000092d_blk00000943 : LUT1
    generic map(
      INIT => X"2"
    )
    port map (
      I0 => sig00000a99,
      O => blk0000092d_sig0000197f
    );
  blk0000092d_blk00000942 : LUT1
    generic map(
      INIT => X"2"
    )
    port map (
      I0 => sig00000a98,
      O => blk0000092d_sig0000197e
    );
  blk0000092d_blk00000941 : LUT1
    generic map(
      INIT => X"2"
    )
    port map (
      I0 => sig00000a97,
      O => blk0000092d_sig0000197d
    );
  blk0000092d_blk00000940 : LUT1
    generic map(
      INIT => X"2"
    )
    port map (
      I0 => sig00000a96,
      O => blk0000092d_sig0000197c
    );
  blk0000092d_blk0000093f : LUT1
    generic map(
      INIT => X"2"
    )
    port map (
      I0 => sig00000a95,
      O => blk0000092d_sig0000197b
    );
  blk0000092d_blk0000093e : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => sig00000aa0,
      D => blk0000092d_sig00001979,
      R => sig000008b6,
      Q => sig00000a87
    );
  blk0000092d_blk0000093d : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => sig00000aa0,
      D => blk0000092d_sig00001974,
      R => sig000008b6,
      Q => sig00000a88
    );
  blk0000092d_blk0000093c : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => sig00000aa0,
      D => blk0000092d_sig00001973,
      R => sig000008b6,
      Q => sig00000a89
    );
  blk0000092d_blk0000093b : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => sig00000aa0,
      D => blk0000092d_sig00001972,
      R => sig000008b6,
      Q => sig00000a8a
    );
  blk0000092d_blk0000093a : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => sig00000aa0,
      D => blk0000092d_sig00001971,
      R => sig000008b6,
      Q => sig00000aa3
    );
  blk0000092d_blk00000939 : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => sig00000aa0,
      D => blk0000092d_sig00001970,
      R => sig000008b6,
      Q => sig00000aa4
    );
  blk0000092d_blk00000938 : MUXCY
    port map (
      CI => sig00000a9b,
      DI => sig00000a99,
      S => blk0000092d_sig0000197f,
      O => blk0000092d_sig0000197a
    );
  blk0000092d_blk00000937 : XORCY
    port map (
      CI => sig00000a9b,
      LI => blk0000092d_sig0000197f,
      O => blk0000092d_sig00001979
    );
  blk0000092d_blk00000936 : MUXCY
    port map (
      CI => blk0000092d_sig0000197a,
      DI => sig00000a98,
      S => blk0000092d_sig0000197e,
      O => blk0000092d_sig00001978
    );
  blk0000092d_blk00000935 : MUXCY
    port map (
      CI => blk0000092d_sig00001978,
      DI => sig00000a97,
      S => blk0000092d_sig0000197d,
      O => blk0000092d_sig00001977
    );
  blk0000092d_blk00000934 : MUXCY
    port map (
      CI => blk0000092d_sig00001977,
      DI => sig00000a96,
      S => blk0000092d_sig0000197c,
      O => blk0000092d_sig00001976
    );
  blk0000092d_blk00000933 : MUXCY
    port map (
      CI => blk0000092d_sig00001976,
      DI => sig00000a95,
      S => blk0000092d_sig0000197b,
      O => blk0000092d_sig00001975
    );
  blk0000092d_blk00000932 : XORCY
    port map (
      CI => blk0000092d_sig0000197a,
      LI => blk0000092d_sig0000197e,
      O => blk0000092d_sig00001974
    );
  blk0000092d_blk00000931 : XORCY
    port map (
      CI => blk0000092d_sig00001978,
      LI => blk0000092d_sig0000197d,
      O => blk0000092d_sig00001973
    );
  blk0000092d_blk00000930 : XORCY
    port map (
      CI => blk0000092d_sig00001977,
      LI => blk0000092d_sig0000197c,
      O => blk0000092d_sig00001972
    );
  blk0000092d_blk0000092f : XORCY
    port map (
      CI => blk0000092d_sig00001976,
      LI => blk0000092d_sig0000197b,
      O => blk0000092d_sig00001971
    );
  blk0000092d_blk0000092e : XORCY
    port map (
      CI => blk0000092d_sig00001975,
      LI => sig00000a94,
      O => blk0000092d_sig00001970
    );
  blk00000955_blk0000096b : LUT1
    generic map(
      INIT => X"2"
    )
    port map (
      I0 => sig00000ab3,
      O => blk00000955_sig0000199f
    );
  blk00000955_blk0000096a : LUT1
    generic map(
      INIT => X"2"
    )
    port map (
      I0 => sig00000ab2,
      O => blk00000955_sig0000199e
    );
  blk00000955_blk00000969 : LUT1
    generic map(
      INIT => X"2"
    )
    port map (
      I0 => sig00000ab1,
      O => blk00000955_sig0000199d
    );
  blk00000955_blk00000968 : LUT1
    generic map(
      INIT => X"2"
    )
    port map (
      I0 => sig00000ab0,
      O => blk00000955_sig0000199c
    );
  blk00000955_blk00000967 : LUT1
    generic map(
      INIT => X"2"
    )
    port map (
      I0 => sig00000aaf,
      O => blk00000955_sig0000199b
    );
  blk00000955_blk00000966 : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => sig00000aba,
      D => blk00000955_sig00001999,
      R => sig000008b6,
      Q => sig00000a82
    );
  blk00000955_blk00000965 : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => sig00000aba,
      D => blk00000955_sig00001994,
      R => sig000008b6,
      Q => sig00000a83
    );
  blk00000955_blk00000964 : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => sig00000aba,
      D => blk00000955_sig00001993,
      R => sig000008b6,
      Q => sig00000a84
    );
  blk00000955_blk00000963 : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => sig00000aba,
      D => blk00000955_sig00001992,
      R => sig000008b6,
      Q => sig00000a85
    );
  blk00000955_blk00000962 : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => sig00000aba,
      D => blk00000955_sig00001991,
      R => sig000008b6,
      Q => sig00000abd
    );
  blk00000955_blk00000961 : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => sig00000aba,
      D => blk00000955_sig00001990,
      R => sig000008b6,
      Q => sig00000abe
    );
  blk00000955_blk00000960 : MUXCY
    port map (
      CI => sig00000ab5,
      DI => sig00000ab3,
      S => blk00000955_sig0000199f,
      O => blk00000955_sig0000199a
    );
  blk00000955_blk0000095f : XORCY
    port map (
      CI => sig00000ab5,
      LI => blk00000955_sig0000199f,
      O => blk00000955_sig00001999
    );
  blk00000955_blk0000095e : MUXCY
    port map (
      CI => blk00000955_sig0000199a,
      DI => sig00000ab2,
      S => blk00000955_sig0000199e,
      O => blk00000955_sig00001998
    );
  blk00000955_blk0000095d : MUXCY
    port map (
      CI => blk00000955_sig00001998,
      DI => sig00000ab1,
      S => blk00000955_sig0000199d,
      O => blk00000955_sig00001997
    );
  blk00000955_blk0000095c : MUXCY
    port map (
      CI => blk00000955_sig00001997,
      DI => sig00000ab0,
      S => blk00000955_sig0000199c,
      O => blk00000955_sig00001996
    );
  blk00000955_blk0000095b : MUXCY
    port map (
      CI => blk00000955_sig00001996,
      DI => sig00000aaf,
      S => blk00000955_sig0000199b,
      O => blk00000955_sig00001995
    );
  blk00000955_blk0000095a : XORCY
    port map (
      CI => blk00000955_sig0000199a,
      LI => blk00000955_sig0000199e,
      O => blk00000955_sig00001994
    );
  blk00000955_blk00000959 : XORCY
    port map (
      CI => blk00000955_sig00001998,
      LI => blk00000955_sig0000199d,
      O => blk00000955_sig00001993
    );
  blk00000955_blk00000958 : XORCY
    port map (
      CI => blk00000955_sig00001997,
      LI => blk00000955_sig0000199c,
      O => blk00000955_sig00001992
    );
  blk00000955_blk00000957 : XORCY
    port map (
      CI => blk00000955_sig00001996,
      LI => blk00000955_sig0000199b,
      O => blk00000955_sig00001991
    );
  blk00000955_blk00000956 : XORCY
    port map (
      CI => blk00000955_sig00001995,
      LI => sig00000aae,
      O => blk00000955_sig00001990
    );
  blk000009b1_blk000009b2_blk000009cc : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk000009b1_blk000009b2_sig000019e2,
      Q => sig00000b3e
    );
  blk000009b1_blk000009b2_blk000009cb : SRLC16E
    generic map(
      INIT => X"0000"
    )
    port map (
      A0 => blk000009b1_blk000009b2_sig000019d5,
      A1 => blk000009b1_blk000009b2_sig000019d6,
      A2 => blk000009b1_blk000009b2_sig000019d6,
      A3 => blk000009b1_blk000009b2_sig000019d5,
      CE => ce,
      CLK => clk,
      D => sig000000f9,
      Q => blk000009b1_blk000009b2_sig000019e2,
      Q15 => NLW_blk000009b1_blk000009b2_blk000009cb_Q15_UNCONNECTED
    );
  blk000009b1_blk000009b2_blk000009ca : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk000009b1_blk000009b2_sig000019e1,
      Q => sig00000b3d
    );
  blk000009b1_blk000009b2_blk000009c9 : SRLC16E
    generic map(
      INIT => X"0000"
    )
    port map (
      A0 => blk000009b1_blk000009b2_sig000019d5,
      A1 => blk000009b1_blk000009b2_sig000019d6,
      A2 => blk000009b1_blk000009b2_sig000019d6,
      A3 => blk000009b1_blk000009b2_sig000019d5,
      CE => ce,
      CLK => clk,
      D => sig000000f8,
      Q => blk000009b1_blk000009b2_sig000019e1,
      Q15 => NLW_blk000009b1_blk000009b2_blk000009c9_Q15_UNCONNECTED
    );
  blk000009b1_blk000009b2_blk000009c8 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk000009b1_blk000009b2_sig000019e0,
      Q => sig00000b3f
    );
  blk000009b1_blk000009b2_blk000009c7 : SRLC16E
    generic map(
      INIT => X"0000"
    )
    port map (
      A0 => blk000009b1_blk000009b2_sig000019d5,
      A1 => blk000009b1_blk000009b2_sig000019d6,
      A2 => blk000009b1_blk000009b2_sig000019d6,
      A3 => blk000009b1_blk000009b2_sig000019d5,
      CE => ce,
      CLK => clk,
      D => sig000000fa,
      Q => blk000009b1_blk000009b2_sig000019e0,
      Q15 => NLW_blk000009b1_blk000009b2_blk000009c7_Q15_UNCONNECTED
    );
  blk000009b1_blk000009b2_blk000009c6 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk000009b1_blk000009b2_sig000019df,
      Q => sig00000b3b
    );
  blk000009b1_blk000009b2_blk000009c5 : SRLC16E
    generic map(
      INIT => X"0000"
    )
    port map (
      A0 => blk000009b1_blk000009b2_sig000019d5,
      A1 => blk000009b1_blk000009b2_sig000019d6,
      A2 => blk000009b1_blk000009b2_sig000019d6,
      A3 => blk000009b1_blk000009b2_sig000019d5,
      CE => ce,
      CLK => clk,
      D => sig000000f6,
      Q => blk000009b1_blk000009b2_sig000019df,
      Q15 => NLW_blk000009b1_blk000009b2_blk000009c5_Q15_UNCONNECTED
    );
  blk000009b1_blk000009b2_blk000009c4 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk000009b1_blk000009b2_sig000019de,
      Q => sig00000b3a
    );
  blk000009b1_blk000009b2_blk000009c3 : SRLC16E
    generic map(
      INIT => X"0000"
    )
    port map (
      A0 => blk000009b1_blk000009b2_sig000019d5,
      A1 => blk000009b1_blk000009b2_sig000019d6,
      A2 => blk000009b1_blk000009b2_sig000019d6,
      A3 => blk000009b1_blk000009b2_sig000019d5,
      CE => ce,
      CLK => clk,
      D => sig000000f5,
      Q => blk000009b1_blk000009b2_sig000019de,
      Q15 => NLW_blk000009b1_blk000009b2_blk000009c3_Q15_UNCONNECTED
    );
  blk000009b1_blk000009b2_blk000009c2 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk000009b1_blk000009b2_sig000019dd,
      Q => sig00000b3c
    );
  blk000009b1_blk000009b2_blk000009c1 : SRLC16E
    generic map(
      INIT => X"0000"
    )
    port map (
      A0 => blk000009b1_blk000009b2_sig000019d5,
      A1 => blk000009b1_blk000009b2_sig000019d6,
      A2 => blk000009b1_blk000009b2_sig000019d6,
      A3 => blk000009b1_blk000009b2_sig000019d5,
      CE => ce,
      CLK => clk,
      D => sig000000f7,
      Q => blk000009b1_blk000009b2_sig000019dd,
      Q15 => NLW_blk000009b1_blk000009b2_blk000009c1_Q15_UNCONNECTED
    );
  blk000009b1_blk000009b2_blk000009c0 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk000009b1_blk000009b2_sig000019dc,
      Q => sig00000b38
    );
  blk000009b1_blk000009b2_blk000009bf : SRLC16E
    generic map(
      INIT => X"0000"
    )
    port map (
      A0 => blk000009b1_blk000009b2_sig000019d5,
      A1 => blk000009b1_blk000009b2_sig000019d6,
      A2 => blk000009b1_blk000009b2_sig000019d6,
      A3 => blk000009b1_blk000009b2_sig000019d5,
      CE => ce,
      CLK => clk,
      D => sig000000f3,
      Q => blk000009b1_blk000009b2_sig000019dc,
      Q15 => NLW_blk000009b1_blk000009b2_blk000009bf_Q15_UNCONNECTED
    );
  blk000009b1_blk000009b2_blk000009be : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk000009b1_blk000009b2_sig000019db,
      Q => sig00000b37
    );
  blk000009b1_blk000009b2_blk000009bd : SRLC16E
    generic map(
      INIT => X"0000"
    )
    port map (
      A0 => blk000009b1_blk000009b2_sig000019d5,
      A1 => blk000009b1_blk000009b2_sig000019d6,
      A2 => blk000009b1_blk000009b2_sig000019d6,
      A3 => blk000009b1_blk000009b2_sig000019d5,
      CE => ce,
      CLK => clk,
      D => sig000000f2,
      Q => blk000009b1_blk000009b2_sig000019db,
      Q15 => NLW_blk000009b1_blk000009b2_blk000009bd_Q15_UNCONNECTED
    );
  blk000009b1_blk000009b2_blk000009bc : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk000009b1_blk000009b2_sig000019da,
      Q => sig00000b39
    );
  blk000009b1_blk000009b2_blk000009bb : SRLC16E
    generic map(
      INIT => X"0000"
    )
    port map (
      A0 => blk000009b1_blk000009b2_sig000019d5,
      A1 => blk000009b1_blk000009b2_sig000019d6,
      A2 => blk000009b1_blk000009b2_sig000019d6,
      A3 => blk000009b1_blk000009b2_sig000019d5,
      CE => ce,
      CLK => clk,
      D => sig000000f4,
      Q => blk000009b1_blk000009b2_sig000019da,
      Q15 => NLW_blk000009b1_blk000009b2_blk000009bb_Q15_UNCONNECTED
    );
  blk000009b1_blk000009b2_blk000009ba : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk000009b1_blk000009b2_sig000019d9,
      Q => sig00000b35
    );
  blk000009b1_blk000009b2_blk000009b9 : SRLC16E
    generic map(
      INIT => X"0000"
    )
    port map (
      A0 => blk000009b1_blk000009b2_sig000019d5,
      A1 => blk000009b1_blk000009b2_sig000019d6,
      A2 => blk000009b1_blk000009b2_sig000019d6,
      A3 => blk000009b1_blk000009b2_sig000019d5,
      CE => ce,
      CLK => clk,
      D => sig000000f0,
      Q => blk000009b1_blk000009b2_sig000019d9,
      Q15 => NLW_blk000009b1_blk000009b2_blk000009b9_Q15_UNCONNECTED
    );
  blk000009b1_blk000009b2_blk000009b8 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk000009b1_blk000009b2_sig000019d8,
      Q => sig00000b34
    );
  blk000009b1_blk000009b2_blk000009b7 : SRLC16E
    generic map(
      INIT => X"0000"
    )
    port map (
      A0 => blk000009b1_blk000009b2_sig000019d5,
      A1 => blk000009b1_blk000009b2_sig000019d6,
      A2 => blk000009b1_blk000009b2_sig000019d6,
      A3 => blk000009b1_blk000009b2_sig000019d5,
      CE => ce,
      CLK => clk,
      D => sig000000ef,
      Q => blk000009b1_blk000009b2_sig000019d8,
      Q15 => NLW_blk000009b1_blk000009b2_blk000009b7_Q15_UNCONNECTED
    );
  blk000009b1_blk000009b2_blk000009b6 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk000009b1_blk000009b2_sig000019d7,
      Q => sig00000b36
    );
  blk000009b1_blk000009b2_blk000009b5 : SRLC16E
    generic map(
      INIT => X"0000"
    )
    port map (
      A0 => blk000009b1_blk000009b2_sig000019d5,
      A1 => blk000009b1_blk000009b2_sig000019d6,
      A2 => blk000009b1_blk000009b2_sig000019d6,
      A3 => blk000009b1_blk000009b2_sig000019d5,
      CE => ce,
      CLK => clk,
      D => sig000000f1,
      Q => blk000009b1_blk000009b2_sig000019d7,
      Q15 => NLW_blk000009b1_blk000009b2_blk000009b5_Q15_UNCONNECTED
    );
  blk000009b1_blk000009b2_blk000009b4 : VCC
    port map (
      P => blk000009b1_blk000009b2_sig000019d6
    );
  blk000009b1_blk000009b2_blk000009b3 : GND
    port map (
      G => blk000009b1_blk000009b2_sig000019d5
    );
  blk000009cd_blk000009ce_blk000009e8 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk000009cd_blk000009ce_sig00001a25,
      Q => sig00000b2f
    );
  blk000009cd_blk000009ce_blk000009e7 : SRLC16E
    generic map(
      INIT => X"0000"
    )
    port map (
      A0 => blk000009cd_blk000009ce_sig00001a18,
      A1 => blk000009cd_blk000009ce_sig00001a19,
      A2 => blk000009cd_blk000009ce_sig00001a19,
      A3 => blk000009cd_blk000009ce_sig00001a18,
      CE => ce,
      CLK => clk,
      D => sig00000b56,
      Q => blk000009cd_blk000009ce_sig00001a25,
      Q15 => NLW_blk000009cd_blk000009ce_blk000009e7_Q15_UNCONNECTED
    );
  blk000009cd_blk000009ce_blk000009e6 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk000009cd_blk000009ce_sig00001a24,
      Q => sig00000b2e
    );
  blk000009cd_blk000009ce_blk000009e5 : SRLC16E
    generic map(
      INIT => X"0000"
    )
    port map (
      A0 => blk000009cd_blk000009ce_sig00001a18,
      A1 => blk000009cd_blk000009ce_sig00001a19,
      A2 => blk000009cd_blk000009ce_sig00001a19,
      A3 => blk000009cd_blk000009ce_sig00001a18,
      CE => ce,
      CLK => clk,
      D => sig00000b55,
      Q => blk000009cd_blk000009ce_sig00001a24,
      Q15 => NLW_blk000009cd_blk000009ce_blk000009e5_Q15_UNCONNECTED
    );
  blk000009cd_blk000009ce_blk000009e4 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk000009cd_blk000009ce_sig00001a23,
      Q => sig00000b30
    );
  blk000009cd_blk000009ce_blk000009e3 : SRLC16E
    generic map(
      INIT => X"0000"
    )
    port map (
      A0 => blk000009cd_blk000009ce_sig00001a18,
      A1 => blk000009cd_blk000009ce_sig00001a19,
      A2 => blk000009cd_blk000009ce_sig00001a19,
      A3 => blk000009cd_blk000009ce_sig00001a18,
      CE => ce,
      CLK => clk,
      D => sig00000b57,
      Q => blk000009cd_blk000009ce_sig00001a23,
      Q15 => NLW_blk000009cd_blk000009ce_blk000009e3_Q15_UNCONNECTED
    );
  blk000009cd_blk000009ce_blk000009e2 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk000009cd_blk000009ce_sig00001a22,
      Q => sig00000b2c
    );
  blk000009cd_blk000009ce_blk000009e1 : SRLC16E
    generic map(
      INIT => X"0000"
    )
    port map (
      A0 => blk000009cd_blk000009ce_sig00001a18,
      A1 => blk000009cd_blk000009ce_sig00001a19,
      A2 => blk000009cd_blk000009ce_sig00001a19,
      A3 => blk000009cd_blk000009ce_sig00001a18,
      CE => ce,
      CLK => clk,
      D => sig00000b53,
      Q => blk000009cd_blk000009ce_sig00001a22,
      Q15 => NLW_blk000009cd_blk000009ce_blk000009e1_Q15_UNCONNECTED
    );
  blk000009cd_blk000009ce_blk000009e0 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk000009cd_blk000009ce_sig00001a21,
      Q => sig00000b2b
    );
  blk000009cd_blk000009ce_blk000009df : SRLC16E
    generic map(
      INIT => X"0000"
    )
    port map (
      A0 => blk000009cd_blk000009ce_sig00001a18,
      A1 => blk000009cd_blk000009ce_sig00001a19,
      A2 => blk000009cd_blk000009ce_sig00001a19,
      A3 => blk000009cd_blk000009ce_sig00001a18,
      CE => ce,
      CLK => clk,
      D => sig00000b52,
      Q => blk000009cd_blk000009ce_sig00001a21,
      Q15 => NLW_blk000009cd_blk000009ce_blk000009df_Q15_UNCONNECTED
    );
  blk000009cd_blk000009ce_blk000009de : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk000009cd_blk000009ce_sig00001a20,
      Q => sig00000b2d
    );
  blk000009cd_blk000009ce_blk000009dd : SRLC16E
    generic map(
      INIT => X"0000"
    )
    port map (
      A0 => blk000009cd_blk000009ce_sig00001a18,
      A1 => blk000009cd_blk000009ce_sig00001a19,
      A2 => blk000009cd_blk000009ce_sig00001a19,
      A3 => blk000009cd_blk000009ce_sig00001a18,
      CE => ce,
      CLK => clk,
      D => sig00000b54,
      Q => blk000009cd_blk000009ce_sig00001a20,
      Q15 => NLW_blk000009cd_blk000009ce_blk000009dd_Q15_UNCONNECTED
    );
  blk000009cd_blk000009ce_blk000009dc : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk000009cd_blk000009ce_sig00001a1f,
      Q => sig00000b29
    );
  blk000009cd_blk000009ce_blk000009db : SRLC16E
    generic map(
      INIT => X"0000"
    )
    port map (
      A0 => blk000009cd_blk000009ce_sig00001a18,
      A1 => blk000009cd_blk000009ce_sig00001a19,
      A2 => blk000009cd_blk000009ce_sig00001a19,
      A3 => blk000009cd_blk000009ce_sig00001a18,
      CE => ce,
      CLK => clk,
      D => sig00000b50,
      Q => blk000009cd_blk000009ce_sig00001a1f,
      Q15 => NLW_blk000009cd_blk000009ce_blk000009db_Q15_UNCONNECTED
    );
  blk000009cd_blk000009ce_blk000009da : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk000009cd_blk000009ce_sig00001a1e,
      Q => sig00000b28
    );
  blk000009cd_blk000009ce_blk000009d9 : SRLC16E
    generic map(
      INIT => X"0000"
    )
    port map (
      A0 => blk000009cd_blk000009ce_sig00001a18,
      A1 => blk000009cd_blk000009ce_sig00001a19,
      A2 => blk000009cd_blk000009ce_sig00001a19,
      A3 => blk000009cd_blk000009ce_sig00001a18,
      CE => ce,
      CLK => clk,
      D => sig00000b4f,
      Q => blk000009cd_blk000009ce_sig00001a1e,
      Q15 => NLW_blk000009cd_blk000009ce_blk000009d9_Q15_UNCONNECTED
    );
  blk000009cd_blk000009ce_blk000009d8 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk000009cd_blk000009ce_sig00001a1d,
      Q => sig00000b2a
    );
  blk000009cd_blk000009ce_blk000009d7 : SRLC16E
    generic map(
      INIT => X"0000"
    )
    port map (
      A0 => blk000009cd_blk000009ce_sig00001a18,
      A1 => blk000009cd_blk000009ce_sig00001a19,
      A2 => blk000009cd_blk000009ce_sig00001a19,
      A3 => blk000009cd_blk000009ce_sig00001a18,
      CE => ce,
      CLK => clk,
      D => sig00000b51,
      Q => blk000009cd_blk000009ce_sig00001a1d,
      Q15 => NLW_blk000009cd_blk000009ce_blk000009d7_Q15_UNCONNECTED
    );
  blk000009cd_blk000009ce_blk000009d6 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk000009cd_blk000009ce_sig00001a1c,
      Q => sig00000b26
    );
  blk000009cd_blk000009ce_blk000009d5 : SRLC16E
    generic map(
      INIT => X"0000"
    )
    port map (
      A0 => blk000009cd_blk000009ce_sig00001a18,
      A1 => blk000009cd_blk000009ce_sig00001a19,
      A2 => blk000009cd_blk000009ce_sig00001a19,
      A3 => blk000009cd_blk000009ce_sig00001a18,
      CE => ce,
      CLK => clk,
      D => sig00000b4d,
      Q => blk000009cd_blk000009ce_sig00001a1c,
      Q15 => NLW_blk000009cd_blk000009ce_blk000009d5_Q15_UNCONNECTED
    );
  blk000009cd_blk000009ce_blk000009d4 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk000009cd_blk000009ce_sig00001a1b,
      Q => sig00000b25
    );
  blk000009cd_blk000009ce_blk000009d3 : SRLC16E
    generic map(
      INIT => X"0000"
    )
    port map (
      A0 => blk000009cd_blk000009ce_sig00001a18,
      A1 => blk000009cd_blk000009ce_sig00001a19,
      A2 => blk000009cd_blk000009ce_sig00001a19,
      A3 => blk000009cd_blk000009ce_sig00001a18,
      CE => ce,
      CLK => clk,
      D => sig00000b4c,
      Q => blk000009cd_blk000009ce_sig00001a1b,
      Q15 => NLW_blk000009cd_blk000009ce_blk000009d3_Q15_UNCONNECTED
    );
  blk000009cd_blk000009ce_blk000009d2 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk000009cd_blk000009ce_sig00001a1a,
      Q => sig00000b27
    );
  blk000009cd_blk000009ce_blk000009d1 : SRLC16E
    generic map(
      INIT => X"0000"
    )
    port map (
      A0 => blk000009cd_blk000009ce_sig00001a18,
      A1 => blk000009cd_blk000009ce_sig00001a19,
      A2 => blk000009cd_blk000009ce_sig00001a19,
      A3 => blk000009cd_blk000009ce_sig00001a18,
      CE => ce,
      CLK => clk,
      D => sig00000b4e,
      Q => blk000009cd_blk000009ce_sig00001a1a,
      Q15 => NLW_blk000009cd_blk000009ce_blk000009d1_Q15_UNCONNECTED
    );
  blk000009cd_blk000009ce_blk000009d0 : VCC
    port map (
      P => blk000009cd_blk000009ce_sig00001a19
    );
  blk000009cd_blk000009ce_blk000009cf : GND
    port map (
      G => blk000009cd_blk000009ce_sig00001a18
    );
  blk000009e9_blk000009ea_blk000009ee : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk000009e9_blk000009ea_sig00001a30,
      Q => sig00000b31
    );
  blk000009e9_blk000009ea_blk000009ed : SRLC16E
    generic map(
      INIT => X"0000"
    )
    port map (
      A0 => blk000009e9_blk000009ea_sig00001a2e,
      A1 => blk000009e9_blk000009ea_sig00001a2f,
      A2 => blk000009e9_blk000009ea_sig00001a2f,
      A3 => blk000009e9_blk000009ea_sig00001a2e,
      CE => ce,
      CLK => clk,
      D => sig00000b32,
      Q => blk000009e9_blk000009ea_sig00001a30,
      Q15 => NLW_blk000009e9_blk000009ea_blk000009ed_Q15_UNCONNECTED
    );
  blk000009e9_blk000009ea_blk000009ec : VCC
    port map (
      P => blk000009e9_blk000009ea_sig00001a2f
    );
  blk000009e9_blk000009ea_blk000009eb : GND
    port map (
      G => blk000009e9_blk000009ea_sig00001a2e
    );
  blk000009ef_blk00000a23 : LUT2
    generic map(
      INIT => X"6"
    )
    port map (
      I0 => sig00000b30,
      I1 => sig00000b4b,
      O => blk000009ef_sig00001a7e
    );
  blk000009ef_blk00000a22 : LUT2
    generic map(
      INIT => X"6"
    )
    port map (
      I0 => sig00000b2e,
      I1 => sig00000b49,
      O => blk000009ef_sig00001a68
    );
  blk000009ef_blk00000a21 : LUT2
    generic map(
      INIT => X"6"
    )
    port map (
      I0 => sig00000b2d,
      I1 => sig00000b48,
      O => blk000009ef_sig00001a69
    );
  blk000009ef_blk00000a20 : LUT2
    generic map(
      INIT => X"6"
    )
    port map (
      I0 => sig00000b2c,
      I1 => sig00000b47,
      O => blk000009ef_sig00001a6a
    );
  blk000009ef_blk00000a1f : LUT2
    generic map(
      INIT => X"6"
    )
    port map (
      I0 => sig00000b2b,
      I1 => sig00000b46,
      O => blk000009ef_sig00001a6b
    );
  blk000009ef_blk00000a1e : LUT2
    generic map(
      INIT => X"6"
    )
    port map (
      I0 => sig00000b2a,
      I1 => sig00000b45,
      O => blk000009ef_sig00001a6c
    );
  blk000009ef_blk00000a1d : LUT2
    generic map(
      INIT => X"6"
    )
    port map (
      I0 => sig00000b29,
      I1 => sig00000b44,
      O => blk000009ef_sig00001a6d
    );
  blk000009ef_blk00000a1c : LUT2
    generic map(
      INIT => X"6"
    )
    port map (
      I0 => sig00000b28,
      I1 => sig00000b43,
      O => blk000009ef_sig00001a6e
    );
  blk000009ef_blk00000a1b : LUT2
    generic map(
      INIT => X"6"
    )
    port map (
      I0 => sig00000b27,
      I1 => sig00000b42,
      O => blk000009ef_sig00001a6f
    );
  blk000009ef_blk00000a1a : LUT2
    generic map(
      INIT => X"6"
    )
    port map (
      I0 => sig00000b26,
      I1 => sig00000b41,
      O => blk000009ef_sig00001a70
    );
  blk000009ef_blk00000a19 : LUT2
    generic map(
      INIT => X"6"
    )
    port map (
      I0 => sig00000b30,
      I1 => sig00000b4b,
      O => blk000009ef_sig00001a66
    );
  blk000009ef_blk00000a18 : LUT2
    generic map(
      INIT => X"6"
    )
    port map (
      I0 => sig00000b2f,
      I1 => sig00000b4a,
      O => blk000009ef_sig00001a67
    );
  blk000009ef_blk00000a17 : LUT2
    generic map(
      INIT => X"6"
    )
    port map (
      I0 => sig00000b25,
      I1 => sig00000b40,
      O => blk000009ef_sig00001a71
    );
  blk000009ef_blk00000a16 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk000009ef_sig00001a65,
      Q => sig00000b18
    );
  blk000009ef_blk00000a15 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk000009ef_sig00001a64,
      Q => sig00000b19
    );
  blk000009ef_blk00000a14 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk000009ef_sig00001a63,
      Q => sig00000b1a
    );
  blk000009ef_blk00000a13 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk000009ef_sig00001a62,
      Q => sig00000b1b
    );
  blk000009ef_blk00000a12 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk000009ef_sig00001a61,
      Q => sig00000b1c
    );
  blk000009ef_blk00000a11 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk000009ef_sig00001a60,
      Q => sig00000b1d
    );
  blk000009ef_blk00000a10 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk000009ef_sig00001a5f,
      Q => sig00000b1e
    );
  blk000009ef_blk00000a0f : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk000009ef_sig00001a5e,
      Q => sig00000b1f
    );
  blk000009ef_blk00000a0e : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk000009ef_sig00001a5d,
      Q => sig00000b20
    );
  blk000009ef_blk00000a0d : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk000009ef_sig00001a5c,
      Q => sig00000b21
    );
  blk000009ef_blk00000a0c : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk000009ef_sig00001a5b,
      Q => sig00000b22
    );
  blk000009ef_blk00000a0b : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk000009ef_sig00001a5a,
      Q => sig00000b23
    );
  blk000009ef_blk00000a0a : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk000009ef_sig00001a59,
      Q => sig00000b24
    );
  blk000009ef_blk00000a09 : MUXCY
    port map (
      CI => blk000009ef_sig00001a58,
      DI => sig00000b25,
      S => blk000009ef_sig00001a71,
      O => blk000009ef_sig00001a7d
    );
  blk000009ef_blk00000a08 : MUXCY
    port map (
      CI => blk000009ef_sig00001a7d,
      DI => sig00000b26,
      S => blk000009ef_sig00001a70,
      O => blk000009ef_sig00001a7c
    );
  blk000009ef_blk00000a07 : MUXCY
    port map (
      CI => blk000009ef_sig00001a7c,
      DI => sig00000b27,
      S => blk000009ef_sig00001a6f,
      O => blk000009ef_sig00001a7b
    );
  blk000009ef_blk00000a06 : MUXCY
    port map (
      CI => blk000009ef_sig00001a7b,
      DI => sig00000b28,
      S => blk000009ef_sig00001a6e,
      O => blk000009ef_sig00001a7a
    );
  blk000009ef_blk00000a05 : MUXCY
    port map (
      CI => blk000009ef_sig00001a7a,
      DI => sig00000b29,
      S => blk000009ef_sig00001a6d,
      O => blk000009ef_sig00001a79
    );
  blk000009ef_blk00000a04 : MUXCY
    port map (
      CI => blk000009ef_sig00001a79,
      DI => sig00000b2a,
      S => blk000009ef_sig00001a6c,
      O => blk000009ef_sig00001a78
    );
  blk000009ef_blk00000a03 : MUXCY
    port map (
      CI => blk000009ef_sig00001a78,
      DI => sig00000b2b,
      S => blk000009ef_sig00001a6b,
      O => blk000009ef_sig00001a77
    );
  blk000009ef_blk00000a02 : MUXCY
    port map (
      CI => blk000009ef_sig00001a77,
      DI => sig00000b2c,
      S => blk000009ef_sig00001a6a,
      O => blk000009ef_sig00001a76
    );
  blk000009ef_blk00000a01 : MUXCY
    port map (
      CI => blk000009ef_sig00001a76,
      DI => sig00000b2d,
      S => blk000009ef_sig00001a69,
      O => blk000009ef_sig00001a75
    );
  blk000009ef_blk00000a00 : MUXCY
    port map (
      CI => blk000009ef_sig00001a75,
      DI => sig00000b2e,
      S => blk000009ef_sig00001a68,
      O => blk000009ef_sig00001a74
    );
  blk000009ef_blk000009ff : MUXCY
    port map (
      CI => blk000009ef_sig00001a74,
      DI => sig00000b2f,
      S => blk000009ef_sig00001a67,
      O => blk000009ef_sig00001a73
    );
  blk000009ef_blk000009fe : MUXCY
    port map (
      CI => blk000009ef_sig00001a73,
      DI => sig00000b30,
      S => blk000009ef_sig00001a7e,
      O => blk000009ef_sig00001a72
    );
  blk000009ef_blk000009fd : XORCY
    port map (
      CI => blk000009ef_sig00001a58,
      LI => blk000009ef_sig00001a71,
      O => blk000009ef_sig00001a65
    );
  blk000009ef_blk000009fc : XORCY
    port map (
      CI => blk000009ef_sig00001a7d,
      LI => blk000009ef_sig00001a70,
      O => blk000009ef_sig00001a64
    );
  blk000009ef_blk000009fb : XORCY
    port map (
      CI => blk000009ef_sig00001a7c,
      LI => blk000009ef_sig00001a6f,
      O => blk000009ef_sig00001a63
    );
  blk000009ef_blk000009fa : XORCY
    port map (
      CI => blk000009ef_sig00001a7b,
      LI => blk000009ef_sig00001a6e,
      O => blk000009ef_sig00001a62
    );
  blk000009ef_blk000009f9 : XORCY
    port map (
      CI => blk000009ef_sig00001a7a,
      LI => blk000009ef_sig00001a6d,
      O => blk000009ef_sig00001a61
    );
  blk000009ef_blk000009f8 : XORCY
    port map (
      CI => blk000009ef_sig00001a79,
      LI => blk000009ef_sig00001a6c,
      O => blk000009ef_sig00001a60
    );
  blk000009ef_blk000009f7 : XORCY
    port map (
      CI => blk000009ef_sig00001a78,
      LI => blk000009ef_sig00001a6b,
      O => blk000009ef_sig00001a5f
    );
  blk000009ef_blk000009f6 : XORCY
    port map (
      CI => blk000009ef_sig00001a77,
      LI => blk000009ef_sig00001a6a,
      O => blk000009ef_sig00001a5e
    );
  blk000009ef_blk000009f5 : XORCY
    port map (
      CI => blk000009ef_sig00001a76,
      LI => blk000009ef_sig00001a69,
      O => blk000009ef_sig00001a5d
    );
  blk000009ef_blk000009f4 : XORCY
    port map (
      CI => blk000009ef_sig00001a75,
      LI => blk000009ef_sig00001a68,
      O => blk000009ef_sig00001a5c
    );
  blk000009ef_blk000009f3 : XORCY
    port map (
      CI => blk000009ef_sig00001a74,
      LI => blk000009ef_sig00001a67,
      O => blk000009ef_sig00001a5b
    );
  blk000009ef_blk000009f2 : XORCY
    port map (
      CI => blk000009ef_sig00001a73,
      LI => blk000009ef_sig00001a7e,
      O => blk000009ef_sig00001a5a
    );
  blk000009ef_blk000009f1 : XORCY
    port map (
      CI => blk000009ef_sig00001a72,
      LI => blk000009ef_sig00001a66,
      O => blk000009ef_sig00001a59
    );
  blk000009ef_blk000009f0 : GND
    port map (
      G => blk000009ef_sig00001a58
    );
  blk00000a24_blk00000a58 : LUT2
    generic map(
      INIT => X"9"
    )
    port map (
      I0 => sig00000b30,
      I1 => sig00000b4b,
      O => blk00000a24_sig00001acc
    );
  blk00000a24_blk00000a57 : LUT2
    generic map(
      INIT => X"9"
    )
    port map (
      I0 => sig00000b2e,
      I1 => sig00000b49,
      O => blk00000a24_sig00001ab5
    );
  blk00000a24_blk00000a56 : LUT2
    generic map(
      INIT => X"9"
    )
    port map (
      I0 => sig00000b2d,
      I1 => sig00000b48,
      O => blk00000a24_sig00001ab6
    );
  blk00000a24_blk00000a55 : LUT2
    generic map(
      INIT => X"9"
    )
    port map (
      I0 => sig00000b2c,
      I1 => sig00000b47,
      O => blk00000a24_sig00001ab7
    );
  blk00000a24_blk00000a54 : LUT2
    generic map(
      INIT => X"9"
    )
    port map (
      I0 => sig00000b2b,
      I1 => sig00000b46,
      O => blk00000a24_sig00001ab8
    );
  blk00000a24_blk00000a53 : LUT2
    generic map(
      INIT => X"9"
    )
    port map (
      I0 => sig00000b2a,
      I1 => sig00000b45,
      O => blk00000a24_sig00001ab9
    );
  blk00000a24_blk00000a52 : LUT2
    generic map(
      INIT => X"9"
    )
    port map (
      I0 => sig00000b29,
      I1 => sig00000b44,
      O => blk00000a24_sig00001aba
    );
  blk00000a24_blk00000a51 : LUT2
    generic map(
      INIT => X"9"
    )
    port map (
      I0 => sig00000b28,
      I1 => sig00000b43,
      O => blk00000a24_sig00001abb
    );
  blk00000a24_blk00000a50 : LUT2
    generic map(
      INIT => X"9"
    )
    port map (
      I0 => sig00000b27,
      I1 => sig00000b42,
      O => blk00000a24_sig00001abc
    );
  blk00000a24_blk00000a4f : LUT2
    generic map(
      INIT => X"9"
    )
    port map (
      I0 => sig00000b26,
      I1 => sig00000b41,
      O => blk00000a24_sig00001abd
    );
  blk00000a24_blk00000a4e : LUT2
    generic map(
      INIT => X"9"
    )
    port map (
      I0 => sig00000b30,
      I1 => sig00000b4b,
      O => blk00000a24_sig00001ab3
    );
  blk00000a24_blk00000a4d : LUT2
    generic map(
      INIT => X"9"
    )
    port map (
      I0 => sig00000b2f,
      I1 => sig00000b4a,
      O => blk00000a24_sig00001ab4
    );
  blk00000a24_blk00000a4c : LUT2
    generic map(
      INIT => X"9"
    )
    port map (
      I0 => sig00000b25,
      I1 => sig00000b40,
      O => blk00000a24_sig00001abe
    );
  blk00000a24_blk00000a4b : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000a24_sig00001ab2,
      Q => sig00000b0b
    );
  blk00000a24_blk00000a4a : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000a24_sig00001ab1,
      Q => sig00000b0c
    );
  blk00000a24_blk00000a49 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000a24_sig00001ab0,
      Q => sig00000b0d
    );
  blk00000a24_blk00000a48 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000a24_sig00001aaf,
      Q => sig00000b0e
    );
  blk00000a24_blk00000a47 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000a24_sig00001aae,
      Q => sig00000b0f
    );
  blk00000a24_blk00000a46 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000a24_sig00001aad,
      Q => sig00000b10
    );
  blk00000a24_blk00000a45 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000a24_sig00001aac,
      Q => sig00000b11
    );
  blk00000a24_blk00000a44 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000a24_sig00001aab,
      Q => sig00000b12
    );
  blk00000a24_blk00000a43 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000a24_sig00001aaa,
      Q => sig00000b13
    );
  blk00000a24_blk00000a42 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000a24_sig00001aa9,
      Q => sig00000b14
    );
  blk00000a24_blk00000a41 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000a24_sig00001aa8,
      Q => sig00000b15
    );
  blk00000a24_blk00000a40 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000a24_sig00001aa7,
      Q => sig00000b16
    );
  blk00000a24_blk00000a3f : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000a24_sig00001aa6,
      Q => sig00000b17
    );
  blk00000a24_blk00000a3e : MUXCY
    port map (
      CI => blk00000a24_sig00001acb,
      DI => sig00000b25,
      S => blk00000a24_sig00001abe,
      O => blk00000a24_sig00001aca
    );
  blk00000a24_blk00000a3d : MUXCY
    port map (
      CI => blk00000a24_sig00001aca,
      DI => sig00000b26,
      S => blk00000a24_sig00001abd,
      O => blk00000a24_sig00001ac9
    );
  blk00000a24_blk00000a3c : MUXCY
    port map (
      CI => blk00000a24_sig00001ac9,
      DI => sig00000b27,
      S => blk00000a24_sig00001abc,
      O => blk00000a24_sig00001ac8
    );
  blk00000a24_blk00000a3b : MUXCY
    port map (
      CI => blk00000a24_sig00001ac8,
      DI => sig00000b28,
      S => blk00000a24_sig00001abb,
      O => blk00000a24_sig00001ac7
    );
  blk00000a24_blk00000a3a : MUXCY
    port map (
      CI => blk00000a24_sig00001ac7,
      DI => sig00000b29,
      S => blk00000a24_sig00001aba,
      O => blk00000a24_sig00001ac6
    );
  blk00000a24_blk00000a39 : MUXCY
    port map (
      CI => blk00000a24_sig00001ac6,
      DI => sig00000b2a,
      S => blk00000a24_sig00001ab9,
      O => blk00000a24_sig00001ac5
    );
  blk00000a24_blk00000a38 : MUXCY
    port map (
      CI => blk00000a24_sig00001ac5,
      DI => sig00000b2b,
      S => blk00000a24_sig00001ab8,
      O => blk00000a24_sig00001ac4
    );
  blk00000a24_blk00000a37 : MUXCY
    port map (
      CI => blk00000a24_sig00001ac4,
      DI => sig00000b2c,
      S => blk00000a24_sig00001ab7,
      O => blk00000a24_sig00001ac3
    );
  blk00000a24_blk00000a36 : MUXCY
    port map (
      CI => blk00000a24_sig00001ac3,
      DI => sig00000b2d,
      S => blk00000a24_sig00001ab6,
      O => blk00000a24_sig00001ac2
    );
  blk00000a24_blk00000a35 : MUXCY
    port map (
      CI => blk00000a24_sig00001ac2,
      DI => sig00000b2e,
      S => blk00000a24_sig00001ab5,
      O => blk00000a24_sig00001ac1
    );
  blk00000a24_blk00000a34 : MUXCY
    port map (
      CI => blk00000a24_sig00001ac1,
      DI => sig00000b2f,
      S => blk00000a24_sig00001ab4,
      O => blk00000a24_sig00001ac0
    );
  blk00000a24_blk00000a33 : MUXCY
    port map (
      CI => blk00000a24_sig00001ac0,
      DI => sig00000b30,
      S => blk00000a24_sig00001acc,
      O => blk00000a24_sig00001abf
    );
  blk00000a24_blk00000a32 : XORCY
    port map (
      CI => blk00000a24_sig00001acb,
      LI => blk00000a24_sig00001abe,
      O => blk00000a24_sig00001ab2
    );
  blk00000a24_blk00000a31 : XORCY
    port map (
      CI => blk00000a24_sig00001aca,
      LI => blk00000a24_sig00001abd,
      O => blk00000a24_sig00001ab1
    );
  blk00000a24_blk00000a30 : XORCY
    port map (
      CI => blk00000a24_sig00001ac9,
      LI => blk00000a24_sig00001abc,
      O => blk00000a24_sig00001ab0
    );
  blk00000a24_blk00000a2f : XORCY
    port map (
      CI => blk00000a24_sig00001ac8,
      LI => blk00000a24_sig00001abb,
      O => blk00000a24_sig00001aaf
    );
  blk00000a24_blk00000a2e : XORCY
    port map (
      CI => blk00000a24_sig00001ac7,
      LI => blk00000a24_sig00001aba,
      O => blk00000a24_sig00001aae
    );
  blk00000a24_blk00000a2d : XORCY
    port map (
      CI => blk00000a24_sig00001ac6,
      LI => blk00000a24_sig00001ab9,
      O => blk00000a24_sig00001aad
    );
  blk00000a24_blk00000a2c : XORCY
    port map (
      CI => blk00000a24_sig00001ac5,
      LI => blk00000a24_sig00001ab8,
      O => blk00000a24_sig00001aac
    );
  blk00000a24_blk00000a2b : XORCY
    port map (
      CI => blk00000a24_sig00001ac4,
      LI => blk00000a24_sig00001ab7,
      O => blk00000a24_sig00001aab
    );
  blk00000a24_blk00000a2a : XORCY
    port map (
      CI => blk00000a24_sig00001ac3,
      LI => blk00000a24_sig00001ab6,
      O => blk00000a24_sig00001aaa
    );
  blk00000a24_blk00000a29 : XORCY
    port map (
      CI => blk00000a24_sig00001ac2,
      LI => blk00000a24_sig00001ab5,
      O => blk00000a24_sig00001aa9
    );
  blk00000a24_blk00000a28 : XORCY
    port map (
      CI => blk00000a24_sig00001ac1,
      LI => blk00000a24_sig00001ab4,
      O => blk00000a24_sig00001aa8
    );
  blk00000a24_blk00000a27 : XORCY
    port map (
      CI => blk00000a24_sig00001ac0,
      LI => blk00000a24_sig00001acc,
      O => blk00000a24_sig00001aa7
    );
  blk00000a24_blk00000a26 : XORCY
    port map (
      CI => blk00000a24_sig00001abf,
      LI => blk00000a24_sig00001ab3,
      O => blk00000a24_sig00001aa6
    );
  blk00000a24_blk00000a25 : VCC
    port map (
      P => blk00000a24_sig00001acb
    );
  blk00000a59_blk00000a5a_blk00000a76 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000a59_blk00000a5a_sig00001b14,
      Q => sig00000b09
    );
  blk00000a59_blk00000a5a_blk00000a75 : SRLC16E
    generic map(
      INIT => X"0000"
    )
    port map (
      A0 => blk00000a59_blk00000a5a_sig00001b06,
      A1 => blk00000a59_blk00000a5a_sig00001b07,
      A2 => blk00000a59_blk00000a5a_sig00001b07,
      A3 => blk00000a59_blk00000a5a_sig00001b06,
      CE => ce,
      CLK => clk,
      D => sig00000b16,
      Q => blk00000a59_blk00000a5a_sig00001b14,
      Q15 => NLW_blk00000a59_blk00000a5a_blk00000a75_Q15_UNCONNECTED
    );
  blk00000a59_blk00000a5a_blk00000a74 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000a59_blk00000a5a_sig00001b13,
      Q => sig00000b08
    );
  blk00000a59_blk00000a5a_blk00000a73 : SRLC16E
    generic map(
      INIT => X"0000"
    )
    port map (
      A0 => blk00000a59_blk00000a5a_sig00001b06,
      A1 => blk00000a59_blk00000a5a_sig00001b07,
      A2 => blk00000a59_blk00000a5a_sig00001b07,
      A3 => blk00000a59_blk00000a5a_sig00001b06,
      CE => ce,
      CLK => clk,
      D => sig00000b15,
      Q => blk00000a59_blk00000a5a_sig00001b13,
      Q15 => NLW_blk00000a59_blk00000a5a_blk00000a73_Q15_UNCONNECTED
    );
  blk00000a59_blk00000a5a_blk00000a72 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000a59_blk00000a5a_sig00001b12,
      Q => sig00000b0a
    );
  blk00000a59_blk00000a5a_blk00000a71 : SRLC16E
    generic map(
      INIT => X"0000"
    )
    port map (
      A0 => blk00000a59_blk00000a5a_sig00001b06,
      A1 => blk00000a59_blk00000a5a_sig00001b07,
      A2 => blk00000a59_blk00000a5a_sig00001b07,
      A3 => blk00000a59_blk00000a5a_sig00001b06,
      CE => ce,
      CLK => clk,
      D => sig00000b17,
      Q => blk00000a59_blk00000a5a_sig00001b12,
      Q15 => NLW_blk00000a59_blk00000a5a_blk00000a71_Q15_UNCONNECTED
    );
  blk00000a59_blk00000a5a_blk00000a70 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000a59_blk00000a5a_sig00001b11,
      Q => sig00000b06
    );
  blk00000a59_blk00000a5a_blk00000a6f : SRLC16E
    generic map(
      INIT => X"0000"
    )
    port map (
      A0 => blk00000a59_blk00000a5a_sig00001b06,
      A1 => blk00000a59_blk00000a5a_sig00001b07,
      A2 => blk00000a59_blk00000a5a_sig00001b07,
      A3 => blk00000a59_blk00000a5a_sig00001b06,
      CE => ce,
      CLK => clk,
      D => sig00000b13,
      Q => blk00000a59_blk00000a5a_sig00001b11,
      Q15 => NLW_blk00000a59_blk00000a5a_blk00000a6f_Q15_UNCONNECTED
    );
  blk00000a59_blk00000a5a_blk00000a6e : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000a59_blk00000a5a_sig00001b10,
      Q => sig00000b05
    );
  blk00000a59_blk00000a5a_blk00000a6d : SRLC16E
    generic map(
      INIT => X"0000"
    )
    port map (
      A0 => blk00000a59_blk00000a5a_sig00001b06,
      A1 => blk00000a59_blk00000a5a_sig00001b07,
      A2 => blk00000a59_blk00000a5a_sig00001b07,
      A3 => blk00000a59_blk00000a5a_sig00001b06,
      CE => ce,
      CLK => clk,
      D => sig00000b12,
      Q => blk00000a59_blk00000a5a_sig00001b10,
      Q15 => NLW_blk00000a59_blk00000a5a_blk00000a6d_Q15_UNCONNECTED
    );
  blk00000a59_blk00000a5a_blk00000a6c : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000a59_blk00000a5a_sig00001b0f,
      Q => sig00000b07
    );
  blk00000a59_blk00000a5a_blk00000a6b : SRLC16E
    generic map(
      INIT => X"0000"
    )
    port map (
      A0 => blk00000a59_blk00000a5a_sig00001b06,
      A1 => blk00000a59_blk00000a5a_sig00001b07,
      A2 => blk00000a59_blk00000a5a_sig00001b07,
      A3 => blk00000a59_blk00000a5a_sig00001b06,
      CE => ce,
      CLK => clk,
      D => sig00000b14,
      Q => blk00000a59_blk00000a5a_sig00001b0f,
      Q15 => NLW_blk00000a59_blk00000a5a_blk00000a6b_Q15_UNCONNECTED
    );
  blk00000a59_blk00000a5a_blk00000a6a : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000a59_blk00000a5a_sig00001b0e,
      Q => sig00000b03
    );
  blk00000a59_blk00000a5a_blk00000a69 : SRLC16E
    generic map(
      INIT => X"0000"
    )
    port map (
      A0 => blk00000a59_blk00000a5a_sig00001b06,
      A1 => blk00000a59_blk00000a5a_sig00001b07,
      A2 => blk00000a59_blk00000a5a_sig00001b07,
      A3 => blk00000a59_blk00000a5a_sig00001b06,
      CE => ce,
      CLK => clk,
      D => sig00000b10,
      Q => blk00000a59_blk00000a5a_sig00001b0e,
      Q15 => NLW_blk00000a59_blk00000a5a_blk00000a69_Q15_UNCONNECTED
    );
  blk00000a59_blk00000a5a_blk00000a68 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000a59_blk00000a5a_sig00001b0d,
      Q => sig00000b02
    );
  blk00000a59_blk00000a5a_blk00000a67 : SRLC16E
    generic map(
      INIT => X"0000"
    )
    port map (
      A0 => blk00000a59_blk00000a5a_sig00001b06,
      A1 => blk00000a59_blk00000a5a_sig00001b07,
      A2 => blk00000a59_blk00000a5a_sig00001b07,
      A3 => blk00000a59_blk00000a5a_sig00001b06,
      CE => ce,
      CLK => clk,
      D => sig00000b0f,
      Q => blk00000a59_blk00000a5a_sig00001b0d,
      Q15 => NLW_blk00000a59_blk00000a5a_blk00000a67_Q15_UNCONNECTED
    );
  blk00000a59_blk00000a5a_blk00000a66 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000a59_blk00000a5a_sig00001b0c,
      Q => sig00000b04
    );
  blk00000a59_blk00000a5a_blk00000a65 : SRLC16E
    generic map(
      INIT => X"0000"
    )
    port map (
      A0 => blk00000a59_blk00000a5a_sig00001b06,
      A1 => blk00000a59_blk00000a5a_sig00001b07,
      A2 => blk00000a59_blk00000a5a_sig00001b07,
      A3 => blk00000a59_blk00000a5a_sig00001b06,
      CE => ce,
      CLK => clk,
      D => sig00000b11,
      Q => blk00000a59_blk00000a5a_sig00001b0c,
      Q15 => NLW_blk00000a59_blk00000a5a_blk00000a65_Q15_UNCONNECTED
    );
  blk00000a59_blk00000a5a_blk00000a64 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000a59_blk00000a5a_sig00001b0b,
      Q => sig00000b01
    );
  blk00000a59_blk00000a5a_blk00000a63 : SRLC16E
    generic map(
      INIT => X"0000"
    )
    port map (
      A0 => blk00000a59_blk00000a5a_sig00001b06,
      A1 => blk00000a59_blk00000a5a_sig00001b07,
      A2 => blk00000a59_blk00000a5a_sig00001b07,
      A3 => blk00000a59_blk00000a5a_sig00001b06,
      CE => ce,
      CLK => clk,
      D => sig00000b0e,
      Q => blk00000a59_blk00000a5a_sig00001b0b,
      Q15 => NLW_blk00000a59_blk00000a5a_blk00000a63_Q15_UNCONNECTED
    );
  blk00000a59_blk00000a5a_blk00000a62 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000a59_blk00000a5a_sig00001b0a,
      Q => sig00000b00
    );
  blk00000a59_blk00000a5a_blk00000a61 : SRLC16E
    generic map(
      INIT => X"0000"
    )
    port map (
      A0 => blk00000a59_blk00000a5a_sig00001b06,
      A1 => blk00000a59_blk00000a5a_sig00001b07,
      A2 => blk00000a59_blk00000a5a_sig00001b07,
      A3 => blk00000a59_blk00000a5a_sig00001b06,
      CE => ce,
      CLK => clk,
      D => sig00000b0d,
      Q => blk00000a59_blk00000a5a_sig00001b0a,
      Q15 => NLW_blk00000a59_blk00000a5a_blk00000a61_Q15_UNCONNECTED
    );
  blk00000a59_blk00000a5a_blk00000a60 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000a59_blk00000a5a_sig00001b09,
      Q => sig00000aff
    );
  blk00000a59_blk00000a5a_blk00000a5f : SRLC16E
    generic map(
      INIT => X"0000"
    )
    port map (
      A0 => blk00000a59_blk00000a5a_sig00001b06,
      A1 => blk00000a59_blk00000a5a_sig00001b07,
      A2 => blk00000a59_blk00000a5a_sig00001b07,
      A3 => blk00000a59_blk00000a5a_sig00001b06,
      CE => ce,
      CLK => clk,
      D => sig00000b0c,
      Q => blk00000a59_blk00000a5a_sig00001b09,
      Q15 => NLW_blk00000a59_blk00000a5a_blk00000a5f_Q15_UNCONNECTED
    );
  blk00000a59_blk00000a5a_blk00000a5e : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000a59_blk00000a5a_sig00001b08,
      Q => sig00000afe
    );
  blk00000a59_blk00000a5a_blk00000a5d : SRLC16E
    generic map(
      INIT => X"0000"
    )
    port map (
      A0 => blk00000a59_blk00000a5a_sig00001b06,
      A1 => blk00000a59_blk00000a5a_sig00001b07,
      A2 => blk00000a59_blk00000a5a_sig00001b07,
      A3 => blk00000a59_blk00000a5a_sig00001b06,
      CE => ce,
      CLK => clk,
      D => sig00000b0b,
      Q => blk00000a59_blk00000a5a_sig00001b08,
      Q15 => NLW_blk00000a59_blk00000a5a_blk00000a5d_Q15_UNCONNECTED
    );
  blk00000a59_blk00000a5a_blk00000a5c : VCC
    port map (
      P => blk00000a59_blk00000a5a_sig00001b07
    );
  blk00000a59_blk00000a5a_blk00000a5b : GND
    port map (
      G => blk00000a59_blk00000a5a_sig00001b06
    );
  blk00000a77_blk00000a78_blk00000a94 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000a77_blk00000a78_sig00001b5c,
      Q => sig00000a7f
    );
  blk00000a77_blk00000a78_blk00000a93 : SRLC16E
    generic map(
      INIT => X"0000"
    )
    port map (
      A0 => blk00000a77_blk00000a78_sig00001b4e,
      A1 => blk00000a77_blk00000a78_sig00001b4f,
      A2 => blk00000a77_blk00000a78_sig00001b4f,
      A3 => blk00000a77_blk00000a78_sig00001b4e,
      CE => ce,
      CLK => clk,
      D => sig00000afc,
      Q => blk00000a77_blk00000a78_sig00001b5c,
      Q15 => NLW_blk00000a77_blk00000a78_blk00000a93_Q15_UNCONNECTED
    );
  blk00000a77_blk00000a78_blk00000a92 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000a77_blk00000a78_sig00001b5b,
      Q => sig00000a7e
    );
  blk00000a77_blk00000a78_blk00000a91 : SRLC16E
    generic map(
      INIT => X"0000"
    )
    port map (
      A0 => blk00000a77_blk00000a78_sig00001b4e,
      A1 => blk00000a77_blk00000a78_sig00001b4f,
      A2 => blk00000a77_blk00000a78_sig00001b4f,
      A3 => blk00000a77_blk00000a78_sig00001b4e,
      CE => ce,
      CLK => clk,
      D => sig00000afb,
      Q => blk00000a77_blk00000a78_sig00001b5b,
      Q15 => NLW_blk00000a77_blk00000a78_blk00000a91_Q15_UNCONNECTED
    );
  blk00000a77_blk00000a78_blk00000a90 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000a77_blk00000a78_sig00001b5a,
      Q => sig00000a80
    );
  blk00000a77_blk00000a78_blk00000a8f : SRLC16E
    generic map(
      INIT => X"0000"
    )
    port map (
      A0 => blk00000a77_blk00000a78_sig00001b4e,
      A1 => blk00000a77_blk00000a78_sig00001b4f,
      A2 => blk00000a77_blk00000a78_sig00001b4f,
      A3 => blk00000a77_blk00000a78_sig00001b4e,
      CE => ce,
      CLK => clk,
      D => sig00000afd,
      Q => blk00000a77_blk00000a78_sig00001b5a,
      Q15 => NLW_blk00000a77_blk00000a78_blk00000a8f_Q15_UNCONNECTED
    );
  blk00000a77_blk00000a78_blk00000a8e : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000a77_blk00000a78_sig00001b59,
      Q => sig00000a7c
    );
  blk00000a77_blk00000a78_blk00000a8d : SRLC16E
    generic map(
      INIT => X"0000"
    )
    port map (
      A0 => blk00000a77_blk00000a78_sig00001b4e,
      A1 => blk00000a77_blk00000a78_sig00001b4f,
      A2 => blk00000a77_blk00000a78_sig00001b4f,
      A3 => blk00000a77_blk00000a78_sig00001b4e,
      CE => ce,
      CLK => clk,
      D => sig00000af9,
      Q => blk00000a77_blk00000a78_sig00001b59,
      Q15 => NLW_blk00000a77_blk00000a78_blk00000a8d_Q15_UNCONNECTED
    );
  blk00000a77_blk00000a78_blk00000a8c : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000a77_blk00000a78_sig00001b58,
      Q => sig00000a7b
    );
  blk00000a77_blk00000a78_blk00000a8b : SRLC16E
    generic map(
      INIT => X"0000"
    )
    port map (
      A0 => blk00000a77_blk00000a78_sig00001b4e,
      A1 => blk00000a77_blk00000a78_sig00001b4f,
      A2 => blk00000a77_blk00000a78_sig00001b4f,
      A3 => blk00000a77_blk00000a78_sig00001b4e,
      CE => ce,
      CLK => clk,
      D => sig00000af8,
      Q => blk00000a77_blk00000a78_sig00001b58,
      Q15 => NLW_blk00000a77_blk00000a78_blk00000a8b_Q15_UNCONNECTED
    );
  blk00000a77_blk00000a78_blk00000a8a : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000a77_blk00000a78_sig00001b57,
      Q => sig00000a7d
    );
  blk00000a77_blk00000a78_blk00000a89 : SRLC16E
    generic map(
      INIT => X"0000"
    )
    port map (
      A0 => blk00000a77_blk00000a78_sig00001b4e,
      A1 => blk00000a77_blk00000a78_sig00001b4f,
      A2 => blk00000a77_blk00000a78_sig00001b4f,
      A3 => blk00000a77_blk00000a78_sig00001b4e,
      CE => ce,
      CLK => clk,
      D => sig00000afa,
      Q => blk00000a77_blk00000a78_sig00001b57,
      Q15 => NLW_blk00000a77_blk00000a78_blk00000a89_Q15_UNCONNECTED
    );
  blk00000a77_blk00000a78_blk00000a88 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000a77_blk00000a78_sig00001b56,
      Q => sig00000a79
    );
  blk00000a77_blk00000a78_blk00000a87 : SRLC16E
    generic map(
      INIT => X"0000"
    )
    port map (
      A0 => blk00000a77_blk00000a78_sig00001b4e,
      A1 => blk00000a77_blk00000a78_sig00001b4f,
      A2 => blk00000a77_blk00000a78_sig00001b4f,
      A3 => blk00000a77_blk00000a78_sig00001b4e,
      CE => ce,
      CLK => clk,
      D => sig00000af6,
      Q => blk00000a77_blk00000a78_sig00001b56,
      Q15 => NLW_blk00000a77_blk00000a78_blk00000a87_Q15_UNCONNECTED
    );
  blk00000a77_blk00000a78_blk00000a86 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000a77_blk00000a78_sig00001b55,
      Q => sig00000a78
    );
  blk00000a77_blk00000a78_blk00000a85 : SRLC16E
    generic map(
      INIT => X"0000"
    )
    port map (
      A0 => blk00000a77_blk00000a78_sig00001b4e,
      A1 => blk00000a77_blk00000a78_sig00001b4f,
      A2 => blk00000a77_blk00000a78_sig00001b4f,
      A3 => blk00000a77_blk00000a78_sig00001b4e,
      CE => ce,
      CLK => clk,
      D => sig00000af5,
      Q => blk00000a77_blk00000a78_sig00001b55,
      Q15 => NLW_blk00000a77_blk00000a78_blk00000a85_Q15_UNCONNECTED
    );
  blk00000a77_blk00000a78_blk00000a84 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000a77_blk00000a78_sig00001b54,
      Q => sig00000a7a
    );
  blk00000a77_blk00000a78_blk00000a83 : SRLC16E
    generic map(
      INIT => X"0000"
    )
    port map (
      A0 => blk00000a77_blk00000a78_sig00001b4e,
      A1 => blk00000a77_blk00000a78_sig00001b4f,
      A2 => blk00000a77_blk00000a78_sig00001b4f,
      A3 => blk00000a77_blk00000a78_sig00001b4e,
      CE => ce,
      CLK => clk,
      D => sig00000af7,
      Q => blk00000a77_blk00000a78_sig00001b54,
      Q15 => NLW_blk00000a77_blk00000a78_blk00000a83_Q15_UNCONNECTED
    );
  blk00000a77_blk00000a78_blk00000a82 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000a77_blk00000a78_sig00001b53,
      Q => sig00000a77
    );
  blk00000a77_blk00000a78_blk00000a81 : SRLC16E
    generic map(
      INIT => X"0000"
    )
    port map (
      A0 => blk00000a77_blk00000a78_sig00001b4e,
      A1 => blk00000a77_blk00000a78_sig00001b4f,
      A2 => blk00000a77_blk00000a78_sig00001b4f,
      A3 => blk00000a77_blk00000a78_sig00001b4e,
      CE => ce,
      CLK => clk,
      D => sig00000af4,
      Q => blk00000a77_blk00000a78_sig00001b53,
      Q15 => NLW_blk00000a77_blk00000a78_blk00000a81_Q15_UNCONNECTED
    );
  blk00000a77_blk00000a78_blk00000a80 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000a77_blk00000a78_sig00001b52,
      Q => sig00000a76
    );
  blk00000a77_blk00000a78_blk00000a7f : SRLC16E
    generic map(
      INIT => X"0000"
    )
    port map (
      A0 => blk00000a77_blk00000a78_sig00001b4e,
      A1 => blk00000a77_blk00000a78_sig00001b4f,
      A2 => blk00000a77_blk00000a78_sig00001b4f,
      A3 => blk00000a77_blk00000a78_sig00001b4e,
      CE => ce,
      CLK => clk,
      D => sig00000af3,
      Q => blk00000a77_blk00000a78_sig00001b52,
      Q15 => NLW_blk00000a77_blk00000a78_blk00000a7f_Q15_UNCONNECTED
    );
  blk00000a77_blk00000a78_blk00000a7e : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000a77_blk00000a78_sig00001b51,
      Q => sig00000a75
    );
  blk00000a77_blk00000a78_blk00000a7d : SRLC16E
    generic map(
      INIT => X"0000"
    )
    port map (
      A0 => blk00000a77_blk00000a78_sig00001b4e,
      A1 => blk00000a77_blk00000a78_sig00001b4f,
      A2 => blk00000a77_blk00000a78_sig00001b4f,
      A3 => blk00000a77_blk00000a78_sig00001b4e,
      CE => ce,
      CLK => clk,
      D => sig00000af2,
      Q => blk00000a77_blk00000a78_sig00001b51,
      Q15 => NLW_blk00000a77_blk00000a78_blk00000a7d_Q15_UNCONNECTED
    );
  blk00000a77_blk00000a78_blk00000a7c : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000a77_blk00000a78_sig00001b50,
      Q => sig00000a74
    );
  blk00000a77_blk00000a78_blk00000a7b : SRLC16E
    generic map(
      INIT => X"0000"
    )
    port map (
      A0 => blk00000a77_blk00000a78_sig00001b4e,
      A1 => blk00000a77_blk00000a78_sig00001b4f,
      A2 => blk00000a77_blk00000a78_sig00001b4f,
      A3 => blk00000a77_blk00000a78_sig00001b4e,
      CE => ce,
      CLK => clk,
      D => sig00000af1,
      Q => blk00000a77_blk00000a78_sig00001b50,
      Q15 => NLW_blk00000a77_blk00000a78_blk00000a7b_Q15_UNCONNECTED
    );
  blk00000a77_blk00000a78_blk00000a7a : VCC
    port map (
      P => blk00000a77_blk00000a78_sig00001b4f
    );
  blk00000a77_blk00000a78_blk00000a79 : GND
    port map (
      G => blk00000a77_blk00000a78_sig00001b4e
    );
  blk00000a95_blk00000a96_blk00000a9c : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000a95_blk00000a96_sig00001b70,
      Q => sig000000ec
    );
  blk00000a95_blk00000a96_blk00000a9b : SRLC32E
    generic map(
      INIT => X"00000000"
    )
    port map (
      CLK => clk,
      D => sig00000a83,
      CE => ce,
      Q => blk00000a95_blk00000a96_sig00001b70,
      Q31 => NLW_blk00000a95_blk00000a96_blk00000a9b_Q31_UNCONNECTED,
      A(4) => blk00000a95_blk00000a96_sig00001b6e,
      A(3) => blk00000a95_blk00000a96_sig00001b6e,
      A(2) => blk00000a95_blk00000a96_sig00001b6d,
      A(1) => blk00000a95_blk00000a96_sig00001b6e,
      A(0) => blk00000a95_blk00000a96_sig00001b6d
    );
  blk00000a95_blk00000a96_blk00000a9a : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000a95_blk00000a96_sig00001b6f,
      Q => sig000000eb
    );
  blk00000a95_blk00000a96_blk00000a99 : SRLC32E
    generic map(
      INIT => X"00000000"
    )
    port map (
      CLK => clk,
      D => sig00000a82,
      CE => ce,
      Q => blk00000a95_blk00000a96_sig00001b6f,
      Q31 => NLW_blk00000a95_blk00000a96_blk00000a99_Q31_UNCONNECTED,
      A(4) => blk00000a95_blk00000a96_sig00001b6e,
      A(3) => blk00000a95_blk00000a96_sig00001b6e,
      A(2) => blk00000a95_blk00000a96_sig00001b6d,
      A(1) => blk00000a95_blk00000a96_sig00001b6e,
      A(0) => blk00000a95_blk00000a96_sig00001b6d
    );
  blk00000a95_blk00000a96_blk00000a98 : VCC
    port map (
      P => blk00000a95_blk00000a96_sig00001b6e
    );
  blk00000a95_blk00000a96_blk00000a97 : GND
    port map (
      G => blk00000a95_blk00000a96_sig00001b6d
    );
  blk00000a9d_blk00000a9e_blk00000aa2 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000a9d_blk00000a9e_sig00001b7b,
      Q => sig000009f5
    );
  blk00000a9d_blk00000a9e_blk00000aa1 : SRLC32E
    generic map(
      INIT => X"00000000"
    )
    port map (
      CLK => clk,
      D => sig00000a81,
      CE => ce,
      Q => blk00000a9d_blk00000a9e_sig00001b7b,
      Q31 => NLW_blk00000a9d_blk00000a9e_blk00000aa1_Q31_UNCONNECTED,
      A(4) => blk00000a9d_blk00000a9e_sig00001b7a,
      A(3) => blk00000a9d_blk00000a9e_sig00001b7a,
      A(2) => blk00000a9d_blk00000a9e_sig00001b79,
      A(1) => blk00000a9d_blk00000a9e_sig00001b79,
      A(0) => blk00000a9d_blk00000a9e_sig00001b7a
    );
  blk00000a9d_blk00000a9e_blk00000aa0 : VCC
    port map (
      P => blk00000a9d_blk00000a9e_sig00001b7a
    );
  blk00000a9d_blk00000a9e_blk00000a9f : GND
    port map (
      G => blk00000a9d_blk00000a9e_sig00001b79
    );
  blk00000aa3_blk00000aa4_blk00000aa8 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000aa3_blk00000aa4_sig00001b86,
      Q => sig00000a5f
    );
  blk00000aa3_blk00000aa4_blk00000aa7 : SRLC16E
    generic map(
      INIT => X"0000"
    )
    port map (
      A0 => blk00000aa3_blk00000aa4_sig00001b85,
      A1 => blk00000aa3_blk00000aa4_sig00001b84,
      A2 => blk00000aa3_blk00000aa4_sig00001b84,
      A3 => blk00000aa3_blk00000aa4_sig00001b85,
      CE => ce,
      CLK => clk,
      D => sig00000a60,
      Q => blk00000aa3_blk00000aa4_sig00001b86,
      Q15 => NLW_blk00000aa3_blk00000aa4_blk00000aa7_Q15_UNCONNECTED
    );
  blk00000aa3_blk00000aa4_blk00000aa6 : VCC
    port map (
      P => blk00000aa3_blk00000aa4_sig00001b85
    );
  blk00000aa3_blk00000aa4_blk00000aa5 : GND
    port map (
      G => blk00000aa3_blk00000aa4_sig00001b84
    );
  blk00000aa9_blk00000aaa_blk00000aae : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000aa9_blk00000aaa_sig00001b91,
      Q => sig000000c9
    );
  blk00000aa9_blk00000aaa_blk00000aad : SRLC32E
    generic map(
      INIT => X"00000000"
    )
    port map (
      CLK => clk,
      D => sig000009f9,
      CE => ce,
      Q => blk00000aa9_blk00000aaa_sig00001b91,
      Q31 => NLW_blk00000aa9_blk00000aaa_blk00000aad_Q31_UNCONNECTED,
      A(4) => blk00000aa9_blk00000aaa_sig00001b90,
      A(3) => blk00000aa9_blk00000aaa_sig00001b90,
      A(2) => blk00000aa9_blk00000aaa_sig00001b8f,
      A(1) => blk00000aa9_blk00000aaa_sig00001b90,
      A(0) => blk00000aa9_blk00000aaa_sig00001b8f
    );
  blk00000aa9_blk00000aaa_blk00000aac : VCC
    port map (
      P => blk00000aa9_blk00000aaa_sig00001b90
    );
  blk00000aa9_blk00000aaa_blk00000aab : GND
    port map (
      G => blk00000aa9_blk00000aaa_sig00001b8f
    );
  blk00000aaf_blk00000ab0_blk00000ab6 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000aaf_blk00000ab0_sig00001ba1,
      Q => sig00000a5a
    );
  blk00000aaf_blk00000ab0_blk00000ab5 : SRLC32E
    generic map(
      INIT => X"00000000"
    )
    port map (
      CLK => clk,
      D => sig00000a5c,
      CE => ce,
      Q => blk00000aaf_blk00000ab0_sig00001ba1,
      Q31 => NLW_blk00000aaf_blk00000ab0_blk00000ab5_Q31_UNCONNECTED,
      A(4) => blk00000aaf_blk00000ab0_sig00001b9f,
      A(3) => blk00000aaf_blk00000ab0_sig00001b9f,
      A(2) => blk00000aaf_blk00000ab0_sig00001b9e,
      A(1) => blk00000aaf_blk00000ab0_sig00001b9e,
      A(0) => blk00000aaf_blk00000ab0_sig00001b9f
    );
  blk00000aaf_blk00000ab0_blk00000ab4 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000aaf_blk00000ab0_sig00001ba0,
      Q => sig00000a59
    );
  blk00000aaf_blk00000ab0_blk00000ab3 : SRLC32E
    generic map(
      INIT => X"00000000"
    )
    port map (
      CLK => clk,
      D => sig00000a5b,
      CE => ce,
      Q => blk00000aaf_blk00000ab0_sig00001ba0,
      Q31 => NLW_blk00000aaf_blk00000ab0_blk00000ab3_Q31_UNCONNECTED,
      A(4) => blk00000aaf_blk00000ab0_sig00001b9f,
      A(3) => blk00000aaf_blk00000ab0_sig00001b9f,
      A(2) => blk00000aaf_blk00000ab0_sig00001b9e,
      A(1) => blk00000aaf_blk00000ab0_sig00001b9e,
      A(0) => blk00000aaf_blk00000ab0_sig00001b9f
    );
  blk00000aaf_blk00000ab0_blk00000ab2 : VCC
    port map (
      P => blk00000aaf_blk00000ab0_sig00001b9f
    );
  blk00000aaf_blk00000ab0_blk00000ab1 : GND
    port map (
      G => blk00000aaf_blk00000ab0_sig00001b9e
    );
  blk00000ab7_blk00000ab8_blk00000abe : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000ab7_blk00000ab8_sig00001bb1,
      Q => sig000000ea
    );
  blk00000ab7_blk00000ab8_blk00000abd : SRLC32E
    generic map(
      INIT => X"00000000"
    )
    port map (
      CLK => clk,
      D => sig00000a5e,
      CE => ce,
      Q => blk00000ab7_blk00000ab8_sig00001bb1,
      Q31 => NLW_blk00000ab7_blk00000ab8_blk00000abd_Q31_UNCONNECTED,
      A(4) => blk00000ab7_blk00000ab8_sig00001baf,
      A(3) => blk00000ab7_blk00000ab8_sig00001baf,
      A(2) => blk00000ab7_blk00000ab8_sig00001bae,
      A(1) => blk00000ab7_blk00000ab8_sig00001baf,
      A(0) => blk00000ab7_blk00000ab8_sig00001bae
    );
  blk00000ab7_blk00000ab8_blk00000abc : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000ab7_blk00000ab8_sig00001bb0,
      Q => sig000000e9
    );
  blk00000ab7_blk00000ab8_blk00000abb : SRLC32E
    generic map(
      INIT => X"00000000"
    )
    port map (
      CLK => clk,
      D => sig00000a5d,
      CE => ce,
      Q => blk00000ab7_blk00000ab8_sig00001bb0,
      Q31 => NLW_blk00000ab7_blk00000ab8_blk00000abb_Q31_UNCONNECTED,
      A(4) => blk00000ab7_blk00000ab8_sig00001baf,
      A(3) => blk00000ab7_blk00000ab8_sig00001baf,
      A(2) => blk00000ab7_blk00000ab8_sig00001bae,
      A(1) => blk00000ab7_blk00000ab8_sig00001baf,
      A(0) => blk00000ab7_blk00000ab8_sig00001bae
    );
  blk00000ab7_blk00000ab8_blk00000aba : VCC
    port map (
      P => blk00000ab7_blk00000ab8_sig00001baf
    );
  blk00000ab7_blk00000ab8_blk00000ab9 : GND
    port map (
      G => blk00000ab7_blk00000ab8_sig00001bae
    );
  blk00000abf_blk00000ac0_blk00000ace : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000abf_blk00000ac0_sig00001bd5,
      Q => sig000000e7
    );
  blk00000abf_blk00000ac0_blk00000acd : SRLC32E
    generic map(
      INIT => X"00000000"
    )
    port map (
      CLK => clk,
      D => sig00000a65,
      CE => ce,
      Q => blk00000abf_blk00000ac0_sig00001bd5,
      Q31 => NLW_blk00000abf_blk00000ac0_blk00000acd_Q31_UNCONNECTED,
      A(4) => blk00000abf_blk00000ac0_sig00001bcf,
      A(3) => blk00000abf_blk00000ac0_sig00001bcf,
      A(2) => blk00000abf_blk00000ac0_sig00001bce,
      A(1) => blk00000abf_blk00000ac0_sig00001bcf,
      A(0) => blk00000abf_blk00000ac0_sig00001bce
    );
  blk00000abf_blk00000ac0_blk00000acc : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000abf_blk00000ac0_sig00001bd4,
      Q => sig000000e6
    );
  blk00000abf_blk00000ac0_blk00000acb : SRLC32E
    generic map(
      INIT => X"00000000"
    )
    port map (
      CLK => clk,
      D => sig00000a64,
      CE => ce,
      Q => blk00000abf_blk00000ac0_sig00001bd4,
      Q31 => NLW_blk00000abf_blk00000ac0_blk00000acb_Q31_UNCONNECTED,
      A(4) => blk00000abf_blk00000ac0_sig00001bcf,
      A(3) => blk00000abf_blk00000ac0_sig00001bcf,
      A(2) => blk00000abf_blk00000ac0_sig00001bce,
      A(1) => blk00000abf_blk00000ac0_sig00001bcf,
      A(0) => blk00000abf_blk00000ac0_sig00001bce
    );
  blk00000abf_blk00000ac0_blk00000aca : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000abf_blk00000ac0_sig00001bd3,
      Q => sig000000e8
    );
  blk00000abf_blk00000ac0_blk00000ac9 : SRLC32E
    generic map(
      INIT => X"00000000"
    )
    port map (
      CLK => clk,
      D => sig00000a66,
      CE => ce,
      Q => blk00000abf_blk00000ac0_sig00001bd3,
      Q31 => NLW_blk00000abf_blk00000ac0_blk00000ac9_Q31_UNCONNECTED,
      A(4) => blk00000abf_blk00000ac0_sig00001bcf,
      A(3) => blk00000abf_blk00000ac0_sig00001bcf,
      A(2) => blk00000abf_blk00000ac0_sig00001bce,
      A(1) => blk00000abf_blk00000ac0_sig00001bcf,
      A(0) => blk00000abf_blk00000ac0_sig00001bce
    );
  blk00000abf_blk00000ac0_blk00000ac8 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000abf_blk00000ac0_sig00001bd2,
      Q => sig000000e4
    );
  blk00000abf_blk00000ac0_blk00000ac7 : SRLC32E
    generic map(
      INIT => X"00000000"
    )
    port map (
      CLK => clk,
      D => sig00000a62,
      CE => ce,
      Q => blk00000abf_blk00000ac0_sig00001bd2,
      Q31 => NLW_blk00000abf_blk00000ac0_blk00000ac7_Q31_UNCONNECTED,
      A(4) => blk00000abf_blk00000ac0_sig00001bcf,
      A(3) => blk00000abf_blk00000ac0_sig00001bcf,
      A(2) => blk00000abf_blk00000ac0_sig00001bce,
      A(1) => blk00000abf_blk00000ac0_sig00001bcf,
      A(0) => blk00000abf_blk00000ac0_sig00001bce
    );
  blk00000abf_blk00000ac0_blk00000ac6 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000abf_blk00000ac0_sig00001bd1,
      Q => sig000000e3
    );
  blk00000abf_blk00000ac0_blk00000ac5 : SRLC32E
    generic map(
      INIT => X"00000000"
    )
    port map (
      CLK => clk,
      D => sig00000a61,
      CE => ce,
      Q => blk00000abf_blk00000ac0_sig00001bd1,
      Q31 => NLW_blk00000abf_blk00000ac0_blk00000ac5_Q31_UNCONNECTED,
      A(4) => blk00000abf_blk00000ac0_sig00001bcf,
      A(3) => blk00000abf_blk00000ac0_sig00001bcf,
      A(2) => blk00000abf_blk00000ac0_sig00001bce,
      A(1) => blk00000abf_blk00000ac0_sig00001bcf,
      A(0) => blk00000abf_blk00000ac0_sig00001bce
    );
  blk00000abf_blk00000ac0_blk00000ac4 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000abf_blk00000ac0_sig00001bd0,
      Q => sig000000e5
    );
  blk00000abf_blk00000ac0_blk00000ac3 : SRLC32E
    generic map(
      INIT => X"00000000"
    )
    port map (
      CLK => clk,
      D => sig00000a63,
      CE => ce,
      Q => blk00000abf_blk00000ac0_sig00001bd0,
      Q31 => NLW_blk00000abf_blk00000ac0_blk00000ac3_Q31_UNCONNECTED,
      A(4) => blk00000abf_blk00000ac0_sig00001bcf,
      A(3) => blk00000abf_blk00000ac0_sig00001bcf,
      A(2) => blk00000abf_blk00000ac0_sig00001bce,
      A(1) => blk00000abf_blk00000ac0_sig00001bcf,
      A(0) => blk00000abf_blk00000ac0_sig00001bce
    );
  blk00000abf_blk00000ac0_blk00000ac2 : VCC
    port map (
      P => blk00000abf_blk00000ac0_sig00001bcf
    );
  blk00000abf_blk00000ac0_blk00000ac1 : GND
    port map (
      G => blk00000abf_blk00000ac0_sig00001bce
    );
  blk00000acf_blk00000ad0_blk00000ad6 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000acf_blk00000ad0_sig00001be9,
      Q => sig00000a58
    );
  blk00000acf_blk00000ad0_blk00000ad5 : SRLC16E
    generic map(
      INIT => X"0000"
    )
    port map (
      A0 => blk00000acf_blk00000ad0_sig00001be6,
      A1 => blk00000acf_blk00000ad0_sig00001be6,
      A2 => blk00000acf_blk00000ad0_sig00001be6,
      A3 => blk00000acf_blk00000ad0_sig00001be7,
      CE => ce,
      CLK => clk,
      D => sig00000a8a,
      Q => blk00000acf_blk00000ad0_sig00001be9,
      Q15 => NLW_blk00000acf_blk00000ad0_blk00000ad5_Q15_UNCONNECTED
    );
  blk00000acf_blk00000ad0_blk00000ad4 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000acf_blk00000ad0_sig00001be8,
      Q => sig00000a57
    );
  blk00000acf_blk00000ad0_blk00000ad3 : SRLC16E
    generic map(
      INIT => X"0000"
    )
    port map (
      A0 => blk00000acf_blk00000ad0_sig00001be6,
      A1 => blk00000acf_blk00000ad0_sig00001be6,
      A2 => blk00000acf_blk00000ad0_sig00001be6,
      A3 => blk00000acf_blk00000ad0_sig00001be7,
      CE => ce,
      CLK => clk,
      D => sig00000a89,
      Q => blk00000acf_blk00000ad0_sig00001be8,
      Q15 => NLW_blk00000acf_blk00000ad0_blk00000ad3_Q15_UNCONNECTED
    );
  blk00000acf_blk00000ad0_blk00000ad2 : VCC
    port map (
      P => blk00000acf_blk00000ad0_sig00001be7
    );
  blk00000acf_blk00000ad0_blk00000ad1 : GND
    port map (
      G => blk00000acf_blk00000ad0_sig00001be6
    );
  blk00000ad7_blk00000b0f : LUT2
    generic map(
      INIT => X"9"
    )
    port map (
      I0 => sig00000c6c,
      I1 => sig00000c42,
      O => blk00000ad7_sig00001c27
    );
  blk00000ad7_blk00000b0e : LUT2
    generic map(
      INIT => X"9"
    )
    port map (
      I0 => sig00000c6b,
      I1 => sig00000c41,
      O => blk00000ad7_sig00001c28
    );
  blk00000ad7_blk00000b0d : LUT2
    generic map(
      INIT => X"9"
    )
    port map (
      I0 => sig00000c6a,
      I1 => sig00000c40,
      O => blk00000ad7_sig00001c29
    );
  blk00000ad7_blk00000b0c : LUT2
    generic map(
      INIT => X"9"
    )
    port map (
      I0 => sig00000c69,
      I1 => sig00000c3f,
      O => blk00000ad7_sig00001c2a
    );
  blk00000ad7_blk00000b0b : LUT2
    generic map(
      INIT => X"9"
    )
    port map (
      I0 => sig00000c68,
      I1 => sig00000c3e,
      O => blk00000ad7_sig00001c2b
    );
  blk00000ad7_blk00000b0a : LUT2
    generic map(
      INIT => X"9"
    )
    port map (
      I0 => sig00000c67,
      I1 => sig00000c3d,
      O => blk00000ad7_sig00001c2c
    );
  blk00000ad7_blk00000b09 : LUT2
    generic map(
      INIT => X"9"
    )
    port map (
      I0 => sig00000c66,
      I1 => sig00000c3c,
      O => blk00000ad7_sig00001c2d
    );
  blk00000ad7_blk00000b08 : LUT2
    generic map(
      INIT => X"9"
    )
    port map (
      I0 => sig00000c65,
      I1 => sig00000c3b,
      O => blk00000ad7_sig00001c2e
    );
  blk00000ad7_blk00000b07 : LUT2
    generic map(
      INIT => X"9"
    )
    port map (
      I0 => sig00000c64,
      I1 => sig00000c3a,
      O => blk00000ad7_sig00001c2f
    );
  blk00000ad7_blk00000b06 : LUT2
    generic map(
      INIT => X"9"
    )
    port map (
      I0 => sig00000c70,
      I1 => sig00000c46,
      O => blk00000ad7_sig00001c30
    );
  blk00000ad7_blk00000b05 : LUT2
    generic map(
      INIT => X"9"
    )
    port map (
      I0 => sig00000c6f,
      I1 => sig00000c45,
      O => blk00000ad7_sig00001c24
    );
  blk00000ad7_blk00000b04 : LUT2
    generic map(
      INIT => X"9"
    )
    port map (
      I0 => sig00000c6e,
      I1 => sig00000c44,
      O => blk00000ad7_sig00001c25
    );
  blk00000ad7_blk00000b03 : LUT2
    generic map(
      INIT => X"9"
    )
    port map (
      I0 => sig00000c6d,
      I1 => sig00000c43,
      O => blk00000ad7_sig00001c26
    );
  blk00000ad7_blk00000b02 : LUT2
    generic map(
      INIT => X"9"
    )
    port map (
      I0 => sig00000c63,
      I1 => sig00000c39,
      O => blk00000ad7_sig00001c31
    );
  blk00000ad7_blk00000b01 : MUXCY
    port map (
      CI => blk00000ad7_sig00001c3f,
      DI => sig00000c63,
      S => blk00000ad7_sig00001c31,
      O => blk00000ad7_sig00001c3e
    );
  blk00000ad7_blk00000b00 : MUXCY
    port map (
      CI => blk00000ad7_sig00001c3e,
      DI => sig00000c64,
      S => blk00000ad7_sig00001c2f,
      O => blk00000ad7_sig00001c3d
    );
  blk00000ad7_blk00000aff : MUXCY
    port map (
      CI => blk00000ad7_sig00001c3d,
      DI => sig00000c65,
      S => blk00000ad7_sig00001c2e,
      O => blk00000ad7_sig00001c3c
    );
  blk00000ad7_blk00000afe : MUXCY
    port map (
      CI => blk00000ad7_sig00001c3c,
      DI => sig00000c66,
      S => blk00000ad7_sig00001c2d,
      O => blk00000ad7_sig00001c3b
    );
  blk00000ad7_blk00000afd : MUXCY
    port map (
      CI => blk00000ad7_sig00001c3b,
      DI => sig00000c67,
      S => blk00000ad7_sig00001c2c,
      O => blk00000ad7_sig00001c3a
    );
  blk00000ad7_blk00000afc : MUXCY
    port map (
      CI => blk00000ad7_sig00001c3a,
      DI => sig00000c68,
      S => blk00000ad7_sig00001c2b,
      O => blk00000ad7_sig00001c39
    );
  blk00000ad7_blk00000afb : MUXCY
    port map (
      CI => blk00000ad7_sig00001c39,
      DI => sig00000c69,
      S => blk00000ad7_sig00001c2a,
      O => blk00000ad7_sig00001c38
    );
  blk00000ad7_blk00000afa : MUXCY
    port map (
      CI => blk00000ad7_sig00001c38,
      DI => sig00000c6a,
      S => blk00000ad7_sig00001c29,
      O => blk00000ad7_sig00001c37
    );
  blk00000ad7_blk00000af9 : MUXCY
    port map (
      CI => blk00000ad7_sig00001c37,
      DI => sig00000c6b,
      S => blk00000ad7_sig00001c28,
      O => blk00000ad7_sig00001c36
    );
  blk00000ad7_blk00000af8 : MUXCY
    port map (
      CI => blk00000ad7_sig00001c36,
      DI => sig00000c6c,
      S => blk00000ad7_sig00001c27,
      O => blk00000ad7_sig00001c35
    );
  blk00000ad7_blk00000af7 : MUXCY
    port map (
      CI => blk00000ad7_sig00001c35,
      DI => sig00000c6d,
      S => blk00000ad7_sig00001c26,
      O => blk00000ad7_sig00001c34
    );
  blk00000ad7_blk00000af6 : MUXCY
    port map (
      CI => blk00000ad7_sig00001c34,
      DI => sig00000c6e,
      S => blk00000ad7_sig00001c25,
      O => blk00000ad7_sig00001c33
    );
  blk00000ad7_blk00000af5 : MUXCY
    port map (
      CI => blk00000ad7_sig00001c33,
      DI => sig00000c6f,
      S => blk00000ad7_sig00001c24,
      O => blk00000ad7_sig00001c32
    );
  blk00000ad7_blk00000af4 : XORCY
    port map (
      CI => blk00000ad7_sig00001c3f,
      LI => blk00000ad7_sig00001c31,
      O => blk00000ad7_sig00001c23
    );
  blk00000ad7_blk00000af3 : XORCY
    port map (
      CI => blk00000ad7_sig00001c3e,
      LI => blk00000ad7_sig00001c2f,
      O => blk00000ad7_sig00001c22
    );
  blk00000ad7_blk00000af2 : XORCY
    port map (
      CI => blk00000ad7_sig00001c3d,
      LI => blk00000ad7_sig00001c2e,
      O => blk00000ad7_sig00001c21
    );
  blk00000ad7_blk00000af1 : XORCY
    port map (
      CI => blk00000ad7_sig00001c3c,
      LI => blk00000ad7_sig00001c2d,
      O => blk00000ad7_sig00001c20
    );
  blk00000ad7_blk00000af0 : XORCY
    port map (
      CI => blk00000ad7_sig00001c3b,
      LI => blk00000ad7_sig00001c2c,
      O => blk00000ad7_sig00001c1f
    );
  blk00000ad7_blk00000aef : XORCY
    port map (
      CI => blk00000ad7_sig00001c3a,
      LI => blk00000ad7_sig00001c2b,
      O => blk00000ad7_sig00001c1e
    );
  blk00000ad7_blk00000aee : XORCY
    port map (
      CI => blk00000ad7_sig00001c39,
      LI => blk00000ad7_sig00001c2a,
      O => blk00000ad7_sig00001c1d
    );
  blk00000ad7_blk00000aed : XORCY
    port map (
      CI => blk00000ad7_sig00001c38,
      LI => blk00000ad7_sig00001c29,
      O => blk00000ad7_sig00001c1c
    );
  blk00000ad7_blk00000aec : XORCY
    port map (
      CI => blk00000ad7_sig00001c37,
      LI => blk00000ad7_sig00001c28,
      O => blk00000ad7_sig00001c1b
    );
  blk00000ad7_blk00000aeb : XORCY
    port map (
      CI => blk00000ad7_sig00001c36,
      LI => blk00000ad7_sig00001c27,
      O => blk00000ad7_sig00001c1a
    );
  blk00000ad7_blk00000aea : XORCY
    port map (
      CI => blk00000ad7_sig00001c35,
      LI => blk00000ad7_sig00001c26,
      O => blk00000ad7_sig00001c19
    );
  blk00000ad7_blk00000ae9 : XORCY
    port map (
      CI => blk00000ad7_sig00001c34,
      LI => blk00000ad7_sig00001c25,
      O => blk00000ad7_sig00001c18
    );
  blk00000ad7_blk00000ae8 : XORCY
    port map (
      CI => blk00000ad7_sig00001c33,
      LI => blk00000ad7_sig00001c24,
      O => blk00000ad7_sig00001c17
    );
  blk00000ad7_blk00000ae7 : XORCY
    port map (
      CI => blk00000ad7_sig00001c32,
      LI => blk00000ad7_sig00001c30,
      O => blk00000ad7_sig00001c16
    );
  blk00000ad7_blk00000ae6 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000ad7_sig00001c16,
      Q => sig00000c2a
    );
  blk00000ad7_blk00000ae5 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000ad7_sig00001c17,
      Q => sig00000c29
    );
  blk00000ad7_blk00000ae4 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000ad7_sig00001c18,
      Q => sig00000c28
    );
  blk00000ad7_blk00000ae3 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000ad7_sig00001c19,
      Q => sig00000c27
    );
  blk00000ad7_blk00000ae2 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000ad7_sig00001c1a,
      Q => sig00000c26
    );
  blk00000ad7_blk00000ae1 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000ad7_sig00001c1b,
      Q => sig00000c25
    );
  blk00000ad7_blk00000ae0 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000ad7_sig00001c1c,
      Q => sig00000c24
    );
  blk00000ad7_blk00000adf : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000ad7_sig00001c1d,
      Q => sig00000c23
    );
  blk00000ad7_blk00000ade : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000ad7_sig00001c1e,
      Q => sig00000c22
    );
  blk00000ad7_blk00000add : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000ad7_sig00001c1f,
      Q => sig00000c21
    );
  blk00000ad7_blk00000adc : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000ad7_sig00001c20,
      Q => sig00000c20
    );
  blk00000ad7_blk00000adb : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000ad7_sig00001c21,
      Q => sig00000c1f
    );
  blk00000ad7_blk00000ada : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000ad7_sig00001c22,
      Q => sig00000c1e
    );
  blk00000ad7_blk00000ad9 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000ad7_sig00001c23,
      Q => sig00000c1d
    );
  blk00000ad7_blk00000ad8 : VCC
    port map (
      P => blk00000ad7_sig00001c3f
    );
  blk00000b10_blk00000b48 : LUT2
    generic map(
      INIT => X"6"
    )
    port map (
      I0 => sig00000c6c,
      I1 => sig00000c42,
      O => blk00000b10_sig00001c7e
    );
  blk00000b10_blk00000b47 : LUT2
    generic map(
      INIT => X"6"
    )
    port map (
      I0 => sig00000c6b,
      I1 => sig00000c41,
      O => blk00000b10_sig00001c7f
    );
  blk00000b10_blk00000b46 : LUT2
    generic map(
      INIT => X"6"
    )
    port map (
      I0 => sig00000c6a,
      I1 => sig00000c40,
      O => blk00000b10_sig00001c80
    );
  blk00000b10_blk00000b45 : LUT2
    generic map(
      INIT => X"6"
    )
    port map (
      I0 => sig00000c69,
      I1 => sig00000c3f,
      O => blk00000b10_sig00001c81
    );
  blk00000b10_blk00000b44 : LUT2
    generic map(
      INIT => X"6"
    )
    port map (
      I0 => sig00000c68,
      I1 => sig00000c3e,
      O => blk00000b10_sig00001c82
    );
  blk00000b10_blk00000b43 : LUT2
    generic map(
      INIT => X"6"
    )
    port map (
      I0 => sig00000c67,
      I1 => sig00000c3d,
      O => blk00000b10_sig00001c83
    );
  blk00000b10_blk00000b42 : LUT2
    generic map(
      INIT => X"6"
    )
    port map (
      I0 => sig00000c66,
      I1 => sig00000c3c,
      O => blk00000b10_sig00001c84
    );
  blk00000b10_blk00000b41 : LUT2
    generic map(
      INIT => X"6"
    )
    port map (
      I0 => sig00000c65,
      I1 => sig00000c3b,
      O => blk00000b10_sig00001c85
    );
  blk00000b10_blk00000b40 : LUT2
    generic map(
      INIT => X"6"
    )
    port map (
      I0 => sig00000c64,
      I1 => sig00000c3a,
      O => blk00000b10_sig00001c86
    );
  blk00000b10_blk00000b3f : LUT2
    generic map(
      INIT => X"6"
    )
    port map (
      I0 => sig00000c70,
      I1 => sig00000c46,
      O => blk00000b10_sig00001c87
    );
  blk00000b10_blk00000b3e : LUT2
    generic map(
      INIT => X"6"
    )
    port map (
      I0 => sig00000c6f,
      I1 => sig00000c45,
      O => blk00000b10_sig00001c7b
    );
  blk00000b10_blk00000b3d : LUT2
    generic map(
      INIT => X"6"
    )
    port map (
      I0 => sig00000c6e,
      I1 => sig00000c44,
      O => blk00000b10_sig00001c7c
    );
  blk00000b10_blk00000b3c : LUT2
    generic map(
      INIT => X"6"
    )
    port map (
      I0 => sig00000c6d,
      I1 => sig00000c43,
      O => blk00000b10_sig00001c7d
    );
  blk00000b10_blk00000b3b : LUT2
    generic map(
      INIT => X"6"
    )
    port map (
      I0 => sig00000c63,
      I1 => sig00000c39,
      O => blk00000b10_sig00001c88
    );
  blk00000b10_blk00000b3a : MUXCY
    port map (
      CI => blk00000b10_sig00001c6c,
      DI => sig00000c63,
      S => blk00000b10_sig00001c88,
      O => blk00000b10_sig00001c95
    );
  blk00000b10_blk00000b39 : MUXCY
    port map (
      CI => blk00000b10_sig00001c95,
      DI => sig00000c64,
      S => blk00000b10_sig00001c86,
      O => blk00000b10_sig00001c94
    );
  blk00000b10_blk00000b38 : MUXCY
    port map (
      CI => blk00000b10_sig00001c94,
      DI => sig00000c65,
      S => blk00000b10_sig00001c85,
      O => blk00000b10_sig00001c93
    );
  blk00000b10_blk00000b37 : MUXCY
    port map (
      CI => blk00000b10_sig00001c93,
      DI => sig00000c66,
      S => blk00000b10_sig00001c84,
      O => blk00000b10_sig00001c92
    );
  blk00000b10_blk00000b36 : MUXCY
    port map (
      CI => blk00000b10_sig00001c92,
      DI => sig00000c67,
      S => blk00000b10_sig00001c83,
      O => blk00000b10_sig00001c91
    );
  blk00000b10_blk00000b35 : MUXCY
    port map (
      CI => blk00000b10_sig00001c91,
      DI => sig00000c68,
      S => blk00000b10_sig00001c82,
      O => blk00000b10_sig00001c90
    );
  blk00000b10_blk00000b34 : MUXCY
    port map (
      CI => blk00000b10_sig00001c90,
      DI => sig00000c69,
      S => blk00000b10_sig00001c81,
      O => blk00000b10_sig00001c8f
    );
  blk00000b10_blk00000b33 : MUXCY
    port map (
      CI => blk00000b10_sig00001c8f,
      DI => sig00000c6a,
      S => blk00000b10_sig00001c80,
      O => blk00000b10_sig00001c8e
    );
  blk00000b10_blk00000b32 : MUXCY
    port map (
      CI => blk00000b10_sig00001c8e,
      DI => sig00000c6b,
      S => blk00000b10_sig00001c7f,
      O => blk00000b10_sig00001c8d
    );
  blk00000b10_blk00000b31 : MUXCY
    port map (
      CI => blk00000b10_sig00001c8d,
      DI => sig00000c6c,
      S => blk00000b10_sig00001c7e,
      O => blk00000b10_sig00001c8c
    );
  blk00000b10_blk00000b30 : MUXCY
    port map (
      CI => blk00000b10_sig00001c8c,
      DI => sig00000c6d,
      S => blk00000b10_sig00001c7d,
      O => blk00000b10_sig00001c8b
    );
  blk00000b10_blk00000b2f : MUXCY
    port map (
      CI => blk00000b10_sig00001c8b,
      DI => sig00000c6e,
      S => blk00000b10_sig00001c7c,
      O => blk00000b10_sig00001c8a
    );
  blk00000b10_blk00000b2e : MUXCY
    port map (
      CI => blk00000b10_sig00001c8a,
      DI => sig00000c6f,
      S => blk00000b10_sig00001c7b,
      O => blk00000b10_sig00001c89
    );
  blk00000b10_blk00000b2d : XORCY
    port map (
      CI => blk00000b10_sig00001c6c,
      LI => blk00000b10_sig00001c88,
      O => blk00000b10_sig00001c7a
    );
  blk00000b10_blk00000b2c : XORCY
    port map (
      CI => blk00000b10_sig00001c95,
      LI => blk00000b10_sig00001c86,
      O => blk00000b10_sig00001c79
    );
  blk00000b10_blk00000b2b : XORCY
    port map (
      CI => blk00000b10_sig00001c94,
      LI => blk00000b10_sig00001c85,
      O => blk00000b10_sig00001c78
    );
  blk00000b10_blk00000b2a : XORCY
    port map (
      CI => blk00000b10_sig00001c93,
      LI => blk00000b10_sig00001c84,
      O => blk00000b10_sig00001c77
    );
  blk00000b10_blk00000b29 : XORCY
    port map (
      CI => blk00000b10_sig00001c92,
      LI => blk00000b10_sig00001c83,
      O => blk00000b10_sig00001c76
    );
  blk00000b10_blk00000b28 : XORCY
    port map (
      CI => blk00000b10_sig00001c91,
      LI => blk00000b10_sig00001c82,
      O => blk00000b10_sig00001c75
    );
  blk00000b10_blk00000b27 : XORCY
    port map (
      CI => blk00000b10_sig00001c90,
      LI => blk00000b10_sig00001c81,
      O => blk00000b10_sig00001c74
    );
  blk00000b10_blk00000b26 : XORCY
    port map (
      CI => blk00000b10_sig00001c8f,
      LI => blk00000b10_sig00001c80,
      O => blk00000b10_sig00001c73
    );
  blk00000b10_blk00000b25 : XORCY
    port map (
      CI => blk00000b10_sig00001c8e,
      LI => blk00000b10_sig00001c7f,
      O => blk00000b10_sig00001c72
    );
  blk00000b10_blk00000b24 : XORCY
    port map (
      CI => blk00000b10_sig00001c8d,
      LI => blk00000b10_sig00001c7e,
      O => blk00000b10_sig00001c71
    );
  blk00000b10_blk00000b23 : XORCY
    port map (
      CI => blk00000b10_sig00001c8c,
      LI => blk00000b10_sig00001c7d,
      O => blk00000b10_sig00001c70
    );
  blk00000b10_blk00000b22 : XORCY
    port map (
      CI => blk00000b10_sig00001c8b,
      LI => blk00000b10_sig00001c7c,
      O => blk00000b10_sig00001c6f
    );
  blk00000b10_blk00000b21 : XORCY
    port map (
      CI => blk00000b10_sig00001c8a,
      LI => blk00000b10_sig00001c7b,
      O => blk00000b10_sig00001c6e
    );
  blk00000b10_blk00000b20 : XORCY
    port map (
      CI => blk00000b10_sig00001c89,
      LI => blk00000b10_sig00001c87,
      O => blk00000b10_sig00001c6d
    );
  blk00000b10_blk00000b1f : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000b10_sig00001c6d,
      Q => sig00000c38
    );
  blk00000b10_blk00000b1e : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000b10_sig00001c6e,
      Q => sig00000c37
    );
  blk00000b10_blk00000b1d : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000b10_sig00001c6f,
      Q => sig00000c36
    );
  blk00000b10_blk00000b1c : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000b10_sig00001c70,
      Q => sig00000c35
    );
  blk00000b10_blk00000b1b : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000b10_sig00001c71,
      Q => sig00000c34
    );
  blk00000b10_blk00000b1a : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000b10_sig00001c72,
      Q => sig00000c33
    );
  blk00000b10_blk00000b19 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000b10_sig00001c73,
      Q => sig00000c32
    );
  blk00000b10_blk00000b18 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000b10_sig00001c74,
      Q => sig00000c31
    );
  blk00000b10_blk00000b17 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000b10_sig00001c75,
      Q => sig00000c30
    );
  blk00000b10_blk00000b16 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000b10_sig00001c76,
      Q => sig00000c2f
    );
  blk00000b10_blk00000b15 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000b10_sig00001c77,
      Q => sig00000c2e
    );
  blk00000b10_blk00000b14 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000b10_sig00001c78,
      Q => sig00000c2d
    );
  blk00000b10_blk00000b13 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000b10_sig00001c79,
      Q => sig00000c2c
    );
  blk00000b10_blk00000b12 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000b10_sig00001c7a,
      Q => sig00000c2b
    );
  blk00000b10_blk00000b11 : GND
    port map (
      G => blk00000b10_sig00001c6c
    );
  blk00000b49_blk00000b4a_blk00000b4d : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000b49_blk00000b4a_sig00001ca6,
      Q => sig00000c8f
    );
  blk00000b49_blk00000b4a_blk00000b4c : SRLC16E
    generic map(
      INIT => X"0000"
    )
    port map (
      A0 => blk00000b49_blk00000b4a_sig00001ca5,
      A1 => blk00000b49_blk00000b4a_sig00001ca5,
      A2 => blk00000b49_blk00000b4a_sig00001ca5,
      A3 => blk00000b49_blk00000b4a_sig00001ca5,
      CE => ce,
      CLK => clk,
      D => sig00000c90,
      Q => blk00000b49_blk00000b4a_sig00001ca6,
      Q15 => NLW_blk00000b49_blk00000b4a_blk00000b4c_Q15_UNCONNECTED
    );
  blk00000b49_blk00000b4a_blk00000b4b : GND
    port map (
      G => blk00000b49_blk00000b4a_sig00001ca5
    );
  blk00000b4e_blk00000b4f_blk00000b52 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000b4e_blk00000b4f_sig00001cb7,
      Q => sig00000c90
    );
  blk00000b4e_blk00000b4f_blk00000b51 : SRLC16E
    generic map(
      INIT => X"0000"
    )
    port map (
      A0 => blk00000b4e_blk00000b4f_sig00001cb6,
      A1 => blk00000b4e_blk00000b4f_sig00001cb6,
      A2 => blk00000b4e_blk00000b4f_sig00001cb6,
      A3 => blk00000b4e_blk00000b4f_sig00001cb6,
      CE => ce,
      CLK => clk,
      D => sig00000c91,
      Q => blk00000b4e_blk00000b4f_sig00001cb7,
      Q15 => NLW_blk00000b4e_blk00000b4f_blk00000b51_Q15_UNCONNECTED
    );
  blk00000b4e_blk00000b4f_blk00000b50 : GND
    port map (
      G => blk00000b4e_blk00000b4f_sig00001cb6
    );
  blk00000b53_blk00000b54_blk00000b58 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000b53_blk00000b54_sig00001cc3,
      Q => sig00000c8e
    );
  blk00000b53_blk00000b54_blk00000b57 : SRLC16E
    generic map(
      INIT => X"0000"
    )
    port map (
      A0 => blk00000b53_blk00000b54_sig00001cc1,
      A1 => blk00000b53_blk00000b54_sig00001cc2,
      A2 => blk00000b53_blk00000b54_sig00001cc1,
      A3 => blk00000b53_blk00000b54_sig00001cc1,
      CE => ce,
      CLK => clk,
      D => sig00000c8f,
      Q => blk00000b53_blk00000b54_sig00001cc3,
      Q15 => NLW_blk00000b53_blk00000b54_blk00000b57_Q15_UNCONNECTED
    );
  blk00000b53_blk00000b54_blk00000b56 : VCC
    port map (
      P => blk00000b53_blk00000b54_sig00001cc2
    );
  blk00000b53_blk00000b54_blk00000b55 : GND
    port map (
      G => blk00000b53_blk00000b54_sig00001cc1
    );
  blk00000c06_blk00000c07_blk00000c25 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000c06_blk00000c07_sig00001d10,
      Q => sig00000c6f
    );
  blk00000c06_blk00000c07_blk00000c24 : SRLC16E
    generic map(
      INIT => X"0000"
    )
    port map (
      A0 => blk00000c06_blk00000c07_sig00001d01,
      A1 => blk00000c06_blk00000c07_sig00001d02,
      A2 => blk00000c06_blk00000c07_sig00001d01,
      A3 => blk00000c06_blk00000c07_sig00001d01,
      CE => ce,
      CLK => clk,
      D => sig00000c53,
      Q => blk00000c06_blk00000c07_sig00001d10,
      Q15 => NLW_blk00000c06_blk00000c07_blk00000c24_Q15_UNCONNECTED
    );
  blk00000c06_blk00000c07_blk00000c23 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000c06_blk00000c07_sig00001d0f,
      Q => sig00000c6e
    );
  blk00000c06_blk00000c07_blk00000c22 : SRLC16E
    generic map(
      INIT => X"0000"
    )
    port map (
      A0 => blk00000c06_blk00000c07_sig00001d01,
      A1 => blk00000c06_blk00000c07_sig00001d02,
      A2 => blk00000c06_blk00000c07_sig00001d01,
      A3 => blk00000c06_blk00000c07_sig00001d01,
      CE => ce,
      CLK => clk,
      D => sig00000c52,
      Q => blk00000c06_blk00000c07_sig00001d0f,
      Q15 => NLW_blk00000c06_blk00000c07_blk00000c22_Q15_UNCONNECTED
    );
  blk00000c06_blk00000c07_blk00000c21 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000c06_blk00000c07_sig00001d0e,
      Q => sig00000c70
    );
  blk00000c06_blk00000c07_blk00000c20 : SRLC16E
    generic map(
      INIT => X"0000"
    )
    port map (
      A0 => blk00000c06_blk00000c07_sig00001d01,
      A1 => blk00000c06_blk00000c07_sig00001d02,
      A2 => blk00000c06_blk00000c07_sig00001d01,
      A3 => blk00000c06_blk00000c07_sig00001d01,
      CE => ce,
      CLK => clk,
      D => sig00000c54,
      Q => blk00000c06_blk00000c07_sig00001d0e,
      Q15 => NLW_blk00000c06_blk00000c07_blk00000c20_Q15_UNCONNECTED
    );
  blk00000c06_blk00000c07_blk00000c1f : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000c06_blk00000c07_sig00001d0d,
      Q => sig00000c6d
    );
  blk00000c06_blk00000c07_blk00000c1e : SRLC16E
    generic map(
      INIT => X"0000"
    )
    port map (
      A0 => blk00000c06_blk00000c07_sig00001d01,
      A1 => blk00000c06_blk00000c07_sig00001d02,
      A2 => blk00000c06_blk00000c07_sig00001d01,
      A3 => blk00000c06_blk00000c07_sig00001d01,
      CE => ce,
      CLK => clk,
      D => sig00000c51,
      Q => blk00000c06_blk00000c07_sig00001d0d,
      Q15 => NLW_blk00000c06_blk00000c07_blk00000c1e_Q15_UNCONNECTED
    );
  blk00000c06_blk00000c07_blk00000c1d : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000c06_blk00000c07_sig00001d0c,
      Q => sig00000c6c
    );
  blk00000c06_blk00000c07_blk00000c1c : SRLC16E
    generic map(
      INIT => X"0000"
    )
    port map (
      A0 => blk00000c06_blk00000c07_sig00001d01,
      A1 => blk00000c06_blk00000c07_sig00001d02,
      A2 => blk00000c06_blk00000c07_sig00001d01,
      A3 => blk00000c06_blk00000c07_sig00001d01,
      CE => ce,
      CLK => clk,
      D => sig00000c50,
      Q => blk00000c06_blk00000c07_sig00001d0c,
      Q15 => NLW_blk00000c06_blk00000c07_blk00000c1c_Q15_UNCONNECTED
    );
  blk00000c06_blk00000c07_blk00000c1b : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000c06_blk00000c07_sig00001d0b,
      Q => sig00000c6b
    );
  blk00000c06_blk00000c07_blk00000c1a : SRLC16E
    generic map(
      INIT => X"0000"
    )
    port map (
      A0 => blk00000c06_blk00000c07_sig00001d01,
      A1 => blk00000c06_blk00000c07_sig00001d02,
      A2 => blk00000c06_blk00000c07_sig00001d01,
      A3 => blk00000c06_blk00000c07_sig00001d01,
      CE => ce,
      CLK => clk,
      D => sig00000c4f,
      Q => blk00000c06_blk00000c07_sig00001d0b,
      Q15 => NLW_blk00000c06_blk00000c07_blk00000c1a_Q15_UNCONNECTED
    );
  blk00000c06_blk00000c07_blk00000c19 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000c06_blk00000c07_sig00001d0a,
      Q => sig00000c6a
    );
  blk00000c06_blk00000c07_blk00000c18 : SRLC16E
    generic map(
      INIT => X"0000"
    )
    port map (
      A0 => blk00000c06_blk00000c07_sig00001d01,
      A1 => blk00000c06_blk00000c07_sig00001d02,
      A2 => blk00000c06_blk00000c07_sig00001d01,
      A3 => blk00000c06_blk00000c07_sig00001d01,
      CE => ce,
      CLK => clk,
      D => sig00000c4e,
      Q => blk00000c06_blk00000c07_sig00001d0a,
      Q15 => NLW_blk00000c06_blk00000c07_blk00000c18_Q15_UNCONNECTED
    );
  blk00000c06_blk00000c07_blk00000c17 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000c06_blk00000c07_sig00001d09,
      Q => sig00000c68
    );
  blk00000c06_blk00000c07_blk00000c16 : SRLC16E
    generic map(
      INIT => X"0000"
    )
    port map (
      A0 => blk00000c06_blk00000c07_sig00001d01,
      A1 => blk00000c06_blk00000c07_sig00001d02,
      A2 => blk00000c06_blk00000c07_sig00001d01,
      A3 => blk00000c06_blk00000c07_sig00001d01,
      CE => ce,
      CLK => clk,
      D => sig00000c4c,
      Q => blk00000c06_blk00000c07_sig00001d09,
      Q15 => NLW_blk00000c06_blk00000c07_blk00000c16_Q15_UNCONNECTED
    );
  blk00000c06_blk00000c07_blk00000c15 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000c06_blk00000c07_sig00001d08,
      Q => sig00000c67
    );
  blk00000c06_blk00000c07_blk00000c14 : SRLC16E
    generic map(
      INIT => X"0000"
    )
    port map (
      A0 => blk00000c06_blk00000c07_sig00001d01,
      A1 => blk00000c06_blk00000c07_sig00001d02,
      A2 => blk00000c06_blk00000c07_sig00001d01,
      A3 => blk00000c06_blk00000c07_sig00001d01,
      CE => ce,
      CLK => clk,
      D => sig00000c4b,
      Q => blk00000c06_blk00000c07_sig00001d08,
      Q15 => NLW_blk00000c06_blk00000c07_blk00000c14_Q15_UNCONNECTED
    );
  blk00000c06_blk00000c07_blk00000c13 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000c06_blk00000c07_sig00001d07,
      Q => sig00000c69
    );
  blk00000c06_blk00000c07_blk00000c12 : SRLC16E
    generic map(
      INIT => X"0000"
    )
    port map (
      A0 => blk00000c06_blk00000c07_sig00001d01,
      A1 => blk00000c06_blk00000c07_sig00001d02,
      A2 => blk00000c06_blk00000c07_sig00001d01,
      A3 => blk00000c06_blk00000c07_sig00001d01,
      CE => ce,
      CLK => clk,
      D => sig00000c4d,
      Q => blk00000c06_blk00000c07_sig00001d07,
      Q15 => NLW_blk00000c06_blk00000c07_blk00000c12_Q15_UNCONNECTED
    );
  blk00000c06_blk00000c07_blk00000c11 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000c06_blk00000c07_sig00001d06,
      Q => sig00000c66
    );
  blk00000c06_blk00000c07_blk00000c10 : SRLC16E
    generic map(
      INIT => X"0000"
    )
    port map (
      A0 => blk00000c06_blk00000c07_sig00001d01,
      A1 => blk00000c06_blk00000c07_sig00001d02,
      A2 => blk00000c06_blk00000c07_sig00001d01,
      A3 => blk00000c06_blk00000c07_sig00001d01,
      CE => ce,
      CLK => clk,
      D => sig00000c4a,
      Q => blk00000c06_blk00000c07_sig00001d06,
      Q15 => NLW_blk00000c06_blk00000c07_blk00000c10_Q15_UNCONNECTED
    );
  blk00000c06_blk00000c07_blk00000c0f : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000c06_blk00000c07_sig00001d05,
      Q => sig00000c65
    );
  blk00000c06_blk00000c07_blk00000c0e : SRLC16E
    generic map(
      INIT => X"0000"
    )
    port map (
      A0 => blk00000c06_blk00000c07_sig00001d01,
      A1 => blk00000c06_blk00000c07_sig00001d02,
      A2 => blk00000c06_blk00000c07_sig00001d01,
      A3 => blk00000c06_blk00000c07_sig00001d01,
      CE => ce,
      CLK => clk,
      D => sig00000c49,
      Q => blk00000c06_blk00000c07_sig00001d05,
      Q15 => NLW_blk00000c06_blk00000c07_blk00000c0e_Q15_UNCONNECTED
    );
  blk00000c06_blk00000c07_blk00000c0d : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000c06_blk00000c07_sig00001d04,
      Q => sig00000c64
    );
  blk00000c06_blk00000c07_blk00000c0c : SRLC16E
    generic map(
      INIT => X"0000"
    )
    port map (
      A0 => blk00000c06_blk00000c07_sig00001d01,
      A1 => blk00000c06_blk00000c07_sig00001d02,
      A2 => blk00000c06_blk00000c07_sig00001d01,
      A3 => blk00000c06_blk00000c07_sig00001d01,
      CE => ce,
      CLK => clk,
      D => sig00000c48,
      Q => blk00000c06_blk00000c07_sig00001d04,
      Q15 => NLW_blk00000c06_blk00000c07_blk00000c0c_Q15_UNCONNECTED
    );
  blk00000c06_blk00000c07_blk00000c0b : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000c06_blk00000c07_sig00001d03,
      Q => sig00000c63
    );
  blk00000c06_blk00000c07_blk00000c0a : SRLC16E
    generic map(
      INIT => X"0000"
    )
    port map (
      A0 => blk00000c06_blk00000c07_sig00001d01,
      A1 => blk00000c06_blk00000c07_sig00001d02,
      A2 => blk00000c06_blk00000c07_sig00001d01,
      A3 => blk00000c06_blk00000c07_sig00001d01,
      CE => ce,
      CLK => clk,
      D => sig00000c47,
      Q => blk00000c06_blk00000c07_sig00001d03,
      Q15 => NLW_blk00000c06_blk00000c07_blk00000c0a_Q15_UNCONNECTED
    );
  blk00000c06_blk00000c07_blk00000c09 : VCC
    port map (
      P => blk00000c06_blk00000c07_sig00001d02
    );
  blk00000c06_blk00000c07_blk00000c08 : GND
    port map (
      G => blk00000c06_blk00000c07_sig00001d01
    );
  blk00000c26_blk00000c27_blk00000c45 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000c26_blk00000c27_sig00001d5d,
      Q => sig00000c61
    );
  blk00000c26_blk00000c27_blk00000c44 : SRLC16E
    generic map(
      INIT => X"0000"
    )
    port map (
      A0 => blk00000c26_blk00000c27_sig00001d4e,
      A1 => blk00000c26_blk00000c27_sig00001d4f,
      A2 => blk00000c26_blk00000c27_sig00001d4e,
      A3 => blk00000c26_blk00000c27_sig00001d4e,
      CE => ce,
      CLK => clk,
      D => sig00000bff,
      Q => blk00000c26_blk00000c27_sig00001d5d,
      Q15 => NLW_blk00000c26_blk00000c27_blk00000c44_Q15_UNCONNECTED
    );
  blk00000c26_blk00000c27_blk00000c43 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000c26_blk00000c27_sig00001d5c,
      Q => sig00000c60
    );
  blk00000c26_blk00000c27_blk00000c42 : SRLC16E
    generic map(
      INIT => X"0000"
    )
    port map (
      A0 => blk00000c26_blk00000c27_sig00001d4e,
      A1 => blk00000c26_blk00000c27_sig00001d4f,
      A2 => blk00000c26_blk00000c27_sig00001d4e,
      A3 => blk00000c26_blk00000c27_sig00001d4e,
      CE => ce,
      CLK => clk,
      D => sig00000bfe,
      Q => blk00000c26_blk00000c27_sig00001d5c,
      Q15 => NLW_blk00000c26_blk00000c27_blk00000c42_Q15_UNCONNECTED
    );
  blk00000c26_blk00000c27_blk00000c41 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000c26_blk00000c27_sig00001d5b,
      Q => sig00000c62
    );
  blk00000c26_blk00000c27_blk00000c40 : SRLC16E
    generic map(
      INIT => X"0000"
    )
    port map (
      A0 => blk00000c26_blk00000c27_sig00001d4e,
      A1 => blk00000c26_blk00000c27_sig00001d4f,
      A2 => blk00000c26_blk00000c27_sig00001d4e,
      A3 => blk00000c26_blk00000c27_sig00001d4e,
      CE => ce,
      CLK => clk,
      D => sig00000c00,
      Q => blk00000c26_blk00000c27_sig00001d5b,
      Q15 => NLW_blk00000c26_blk00000c27_blk00000c40_Q15_UNCONNECTED
    );
  blk00000c26_blk00000c27_blk00000c3f : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000c26_blk00000c27_sig00001d5a,
      Q => sig00000c5f
    );
  blk00000c26_blk00000c27_blk00000c3e : SRLC16E
    generic map(
      INIT => X"0000"
    )
    port map (
      A0 => blk00000c26_blk00000c27_sig00001d4e,
      A1 => blk00000c26_blk00000c27_sig00001d4f,
      A2 => blk00000c26_blk00000c27_sig00001d4e,
      A3 => blk00000c26_blk00000c27_sig00001d4e,
      CE => ce,
      CLK => clk,
      D => sig00000bfd,
      Q => blk00000c26_blk00000c27_sig00001d5a,
      Q15 => NLW_blk00000c26_blk00000c27_blk00000c3e_Q15_UNCONNECTED
    );
  blk00000c26_blk00000c27_blk00000c3d : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000c26_blk00000c27_sig00001d59,
      Q => sig00000c5e
    );
  blk00000c26_blk00000c27_blk00000c3c : SRLC16E
    generic map(
      INIT => X"0000"
    )
    port map (
      A0 => blk00000c26_blk00000c27_sig00001d4e,
      A1 => blk00000c26_blk00000c27_sig00001d4f,
      A2 => blk00000c26_blk00000c27_sig00001d4e,
      A3 => blk00000c26_blk00000c27_sig00001d4e,
      CE => ce,
      CLK => clk,
      D => sig00000bfc,
      Q => blk00000c26_blk00000c27_sig00001d59,
      Q15 => NLW_blk00000c26_blk00000c27_blk00000c3c_Q15_UNCONNECTED
    );
  blk00000c26_blk00000c27_blk00000c3b : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000c26_blk00000c27_sig00001d58,
      Q => sig00000c5d
    );
  blk00000c26_blk00000c27_blk00000c3a : SRLC16E
    generic map(
      INIT => X"0000"
    )
    port map (
      A0 => blk00000c26_blk00000c27_sig00001d4e,
      A1 => blk00000c26_blk00000c27_sig00001d4f,
      A2 => blk00000c26_blk00000c27_sig00001d4e,
      A3 => blk00000c26_blk00000c27_sig00001d4e,
      CE => ce,
      CLK => clk,
      D => sig00000bfb,
      Q => blk00000c26_blk00000c27_sig00001d58,
      Q15 => NLW_blk00000c26_blk00000c27_blk00000c3a_Q15_UNCONNECTED
    );
  blk00000c26_blk00000c27_blk00000c39 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000c26_blk00000c27_sig00001d57,
      Q => sig00000c5c
    );
  blk00000c26_blk00000c27_blk00000c38 : SRLC16E
    generic map(
      INIT => X"0000"
    )
    port map (
      A0 => blk00000c26_blk00000c27_sig00001d4e,
      A1 => blk00000c26_blk00000c27_sig00001d4f,
      A2 => blk00000c26_blk00000c27_sig00001d4e,
      A3 => blk00000c26_blk00000c27_sig00001d4e,
      CE => ce,
      CLK => clk,
      D => sig00000bfa,
      Q => blk00000c26_blk00000c27_sig00001d57,
      Q15 => NLW_blk00000c26_blk00000c27_blk00000c38_Q15_UNCONNECTED
    );
  blk00000c26_blk00000c27_blk00000c37 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000c26_blk00000c27_sig00001d56,
      Q => sig00000c5a
    );
  blk00000c26_blk00000c27_blk00000c36 : SRLC16E
    generic map(
      INIT => X"0000"
    )
    port map (
      A0 => blk00000c26_blk00000c27_sig00001d4e,
      A1 => blk00000c26_blk00000c27_sig00001d4f,
      A2 => blk00000c26_blk00000c27_sig00001d4e,
      A3 => blk00000c26_blk00000c27_sig00001d4e,
      CE => ce,
      CLK => clk,
      D => sig00000bf8,
      Q => blk00000c26_blk00000c27_sig00001d56,
      Q15 => NLW_blk00000c26_blk00000c27_blk00000c36_Q15_UNCONNECTED
    );
  blk00000c26_blk00000c27_blk00000c35 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000c26_blk00000c27_sig00001d55,
      Q => sig00000c59
    );
  blk00000c26_blk00000c27_blk00000c34 : SRLC16E
    generic map(
      INIT => X"0000"
    )
    port map (
      A0 => blk00000c26_blk00000c27_sig00001d4e,
      A1 => blk00000c26_blk00000c27_sig00001d4f,
      A2 => blk00000c26_blk00000c27_sig00001d4e,
      A3 => blk00000c26_blk00000c27_sig00001d4e,
      CE => ce,
      CLK => clk,
      D => sig00000bf7,
      Q => blk00000c26_blk00000c27_sig00001d55,
      Q15 => NLW_blk00000c26_blk00000c27_blk00000c34_Q15_UNCONNECTED
    );
  blk00000c26_blk00000c27_blk00000c33 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000c26_blk00000c27_sig00001d54,
      Q => sig00000c5b
    );
  blk00000c26_blk00000c27_blk00000c32 : SRLC16E
    generic map(
      INIT => X"0000"
    )
    port map (
      A0 => blk00000c26_blk00000c27_sig00001d4e,
      A1 => blk00000c26_blk00000c27_sig00001d4f,
      A2 => blk00000c26_blk00000c27_sig00001d4e,
      A3 => blk00000c26_blk00000c27_sig00001d4e,
      CE => ce,
      CLK => clk,
      D => sig00000bf9,
      Q => blk00000c26_blk00000c27_sig00001d54,
      Q15 => NLW_blk00000c26_blk00000c27_blk00000c32_Q15_UNCONNECTED
    );
  blk00000c26_blk00000c27_blk00000c31 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000c26_blk00000c27_sig00001d53,
      Q => sig00000c58
    );
  blk00000c26_blk00000c27_blk00000c30 : SRLC16E
    generic map(
      INIT => X"0000"
    )
    port map (
      A0 => blk00000c26_blk00000c27_sig00001d4e,
      A1 => blk00000c26_blk00000c27_sig00001d4f,
      A2 => blk00000c26_blk00000c27_sig00001d4e,
      A3 => blk00000c26_blk00000c27_sig00001d4e,
      CE => ce,
      CLK => clk,
      D => sig00000bf6,
      Q => blk00000c26_blk00000c27_sig00001d53,
      Q15 => NLW_blk00000c26_blk00000c27_blk00000c30_Q15_UNCONNECTED
    );
  blk00000c26_blk00000c27_blk00000c2f : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000c26_blk00000c27_sig00001d52,
      Q => sig00000c57
    );
  blk00000c26_blk00000c27_blk00000c2e : SRLC16E
    generic map(
      INIT => X"0000"
    )
    port map (
      A0 => blk00000c26_blk00000c27_sig00001d4e,
      A1 => blk00000c26_blk00000c27_sig00001d4f,
      A2 => blk00000c26_blk00000c27_sig00001d4e,
      A3 => blk00000c26_blk00000c27_sig00001d4e,
      CE => ce,
      CLK => clk,
      D => sig00000bf5,
      Q => blk00000c26_blk00000c27_sig00001d52,
      Q15 => NLW_blk00000c26_blk00000c27_blk00000c2e_Q15_UNCONNECTED
    );
  blk00000c26_blk00000c27_blk00000c2d : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000c26_blk00000c27_sig00001d51,
      Q => sig00000c56
    );
  blk00000c26_blk00000c27_blk00000c2c : SRLC16E
    generic map(
      INIT => X"0000"
    )
    port map (
      A0 => blk00000c26_blk00000c27_sig00001d4e,
      A1 => blk00000c26_blk00000c27_sig00001d4f,
      A2 => blk00000c26_blk00000c27_sig00001d4e,
      A3 => blk00000c26_blk00000c27_sig00001d4e,
      CE => ce,
      CLK => clk,
      D => sig00000bf4,
      Q => blk00000c26_blk00000c27_sig00001d51,
      Q15 => NLW_blk00000c26_blk00000c27_blk00000c2c_Q15_UNCONNECTED
    );
  blk00000c26_blk00000c27_blk00000c2b : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000c26_blk00000c27_sig00001d50,
      Q => sig00000c55
    );
  blk00000c26_blk00000c27_blk00000c2a : SRLC16E
    generic map(
      INIT => X"0000"
    )
    port map (
      A0 => blk00000c26_blk00000c27_sig00001d4e,
      A1 => blk00000c26_blk00000c27_sig00001d4f,
      A2 => blk00000c26_blk00000c27_sig00001d4e,
      A3 => blk00000c26_blk00000c27_sig00001d4e,
      CE => ce,
      CLK => clk,
      D => sig00000bf3,
      Q => blk00000c26_blk00000c27_sig00001d50,
      Q15 => NLW_blk00000c26_blk00000c27_blk00000c2a_Q15_UNCONNECTED
    );
  blk00000c26_blk00000c27_blk00000c29 : VCC
    port map (
      P => blk00000c26_blk00000c27_sig00001d4f
    );
  blk00000c26_blk00000c27_blk00000c28 : GND
    port map (
      G => blk00000c26_blk00000c27_sig00001d4e
    );
  blk00000c46_blk00000c47_blk00000c65 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000c46_blk00000c47_sig00001daa,
      Q => sig00000c1b
    );
  blk00000c46_blk00000c47_blk00000c64 : SRLC16E
    generic map(
      INIT => X"0000"
    )
    port map (
      A0 => blk00000c46_blk00000c47_sig00001d9b,
      A1 => blk00000c46_blk00000c47_sig00001d9c,
      A2 => blk00000c46_blk00000c47_sig00001d9b,
      A3 => blk00000c46_blk00000c47_sig00001d9b,
      CE => ce,
      CLK => clk,
      D => sig00000c29,
      Q => blk00000c46_blk00000c47_sig00001daa,
      Q15 => NLW_blk00000c46_blk00000c47_blk00000c64_Q15_UNCONNECTED
    );
  blk00000c46_blk00000c47_blk00000c63 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000c46_blk00000c47_sig00001da9,
      Q => sig00000c1a
    );
  blk00000c46_blk00000c47_blk00000c62 : SRLC16E
    generic map(
      INIT => X"0000"
    )
    port map (
      A0 => blk00000c46_blk00000c47_sig00001d9b,
      A1 => blk00000c46_blk00000c47_sig00001d9c,
      A2 => blk00000c46_blk00000c47_sig00001d9b,
      A3 => blk00000c46_blk00000c47_sig00001d9b,
      CE => ce,
      CLK => clk,
      D => sig00000c28,
      Q => blk00000c46_blk00000c47_sig00001da9,
      Q15 => NLW_blk00000c46_blk00000c47_blk00000c62_Q15_UNCONNECTED
    );
  blk00000c46_blk00000c47_blk00000c61 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000c46_blk00000c47_sig00001da8,
      Q => sig00000c1c
    );
  blk00000c46_blk00000c47_blk00000c60 : SRLC16E
    generic map(
      INIT => X"0000"
    )
    port map (
      A0 => blk00000c46_blk00000c47_sig00001d9b,
      A1 => blk00000c46_blk00000c47_sig00001d9c,
      A2 => blk00000c46_blk00000c47_sig00001d9b,
      A3 => blk00000c46_blk00000c47_sig00001d9b,
      CE => ce,
      CLK => clk,
      D => sig00000c2a,
      Q => blk00000c46_blk00000c47_sig00001da8,
      Q15 => NLW_blk00000c46_blk00000c47_blk00000c60_Q15_UNCONNECTED
    );
  blk00000c46_blk00000c47_blk00000c5f : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000c46_blk00000c47_sig00001da7,
      Q => sig00000c19
    );
  blk00000c46_blk00000c47_blk00000c5e : SRLC16E
    generic map(
      INIT => X"0000"
    )
    port map (
      A0 => blk00000c46_blk00000c47_sig00001d9b,
      A1 => blk00000c46_blk00000c47_sig00001d9c,
      A2 => blk00000c46_blk00000c47_sig00001d9b,
      A3 => blk00000c46_blk00000c47_sig00001d9b,
      CE => ce,
      CLK => clk,
      D => sig00000c27,
      Q => blk00000c46_blk00000c47_sig00001da7,
      Q15 => NLW_blk00000c46_blk00000c47_blk00000c5e_Q15_UNCONNECTED
    );
  blk00000c46_blk00000c47_blk00000c5d : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000c46_blk00000c47_sig00001da6,
      Q => sig00000c18
    );
  blk00000c46_blk00000c47_blk00000c5c : SRLC16E
    generic map(
      INIT => X"0000"
    )
    port map (
      A0 => blk00000c46_blk00000c47_sig00001d9b,
      A1 => blk00000c46_blk00000c47_sig00001d9c,
      A2 => blk00000c46_blk00000c47_sig00001d9b,
      A3 => blk00000c46_blk00000c47_sig00001d9b,
      CE => ce,
      CLK => clk,
      D => sig00000c26,
      Q => blk00000c46_blk00000c47_sig00001da6,
      Q15 => NLW_blk00000c46_blk00000c47_blk00000c5c_Q15_UNCONNECTED
    );
  blk00000c46_blk00000c47_blk00000c5b : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000c46_blk00000c47_sig00001da5,
      Q => sig00000c17
    );
  blk00000c46_blk00000c47_blk00000c5a : SRLC16E
    generic map(
      INIT => X"0000"
    )
    port map (
      A0 => blk00000c46_blk00000c47_sig00001d9b,
      A1 => blk00000c46_blk00000c47_sig00001d9c,
      A2 => blk00000c46_blk00000c47_sig00001d9b,
      A3 => blk00000c46_blk00000c47_sig00001d9b,
      CE => ce,
      CLK => clk,
      D => sig00000c25,
      Q => blk00000c46_blk00000c47_sig00001da5,
      Q15 => NLW_blk00000c46_blk00000c47_blk00000c5a_Q15_UNCONNECTED
    );
  blk00000c46_blk00000c47_blk00000c59 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000c46_blk00000c47_sig00001da4,
      Q => sig00000c16
    );
  blk00000c46_blk00000c47_blk00000c58 : SRLC16E
    generic map(
      INIT => X"0000"
    )
    port map (
      A0 => blk00000c46_blk00000c47_sig00001d9b,
      A1 => blk00000c46_blk00000c47_sig00001d9c,
      A2 => blk00000c46_blk00000c47_sig00001d9b,
      A3 => blk00000c46_blk00000c47_sig00001d9b,
      CE => ce,
      CLK => clk,
      D => sig00000c24,
      Q => blk00000c46_blk00000c47_sig00001da4,
      Q15 => NLW_blk00000c46_blk00000c47_blk00000c58_Q15_UNCONNECTED
    );
  blk00000c46_blk00000c47_blk00000c57 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000c46_blk00000c47_sig00001da3,
      Q => sig00000c14
    );
  blk00000c46_blk00000c47_blk00000c56 : SRLC16E
    generic map(
      INIT => X"0000"
    )
    port map (
      A0 => blk00000c46_blk00000c47_sig00001d9b,
      A1 => blk00000c46_blk00000c47_sig00001d9c,
      A2 => blk00000c46_blk00000c47_sig00001d9b,
      A3 => blk00000c46_blk00000c47_sig00001d9b,
      CE => ce,
      CLK => clk,
      D => sig00000c22,
      Q => blk00000c46_blk00000c47_sig00001da3,
      Q15 => NLW_blk00000c46_blk00000c47_blk00000c56_Q15_UNCONNECTED
    );
  blk00000c46_blk00000c47_blk00000c55 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000c46_blk00000c47_sig00001da2,
      Q => sig00000c13
    );
  blk00000c46_blk00000c47_blk00000c54 : SRLC16E
    generic map(
      INIT => X"0000"
    )
    port map (
      A0 => blk00000c46_blk00000c47_sig00001d9b,
      A1 => blk00000c46_blk00000c47_sig00001d9c,
      A2 => blk00000c46_blk00000c47_sig00001d9b,
      A3 => blk00000c46_blk00000c47_sig00001d9b,
      CE => ce,
      CLK => clk,
      D => sig00000c21,
      Q => blk00000c46_blk00000c47_sig00001da2,
      Q15 => NLW_blk00000c46_blk00000c47_blk00000c54_Q15_UNCONNECTED
    );
  blk00000c46_blk00000c47_blk00000c53 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000c46_blk00000c47_sig00001da1,
      Q => sig00000c15
    );
  blk00000c46_blk00000c47_blk00000c52 : SRLC16E
    generic map(
      INIT => X"0000"
    )
    port map (
      A0 => blk00000c46_blk00000c47_sig00001d9b,
      A1 => blk00000c46_blk00000c47_sig00001d9c,
      A2 => blk00000c46_blk00000c47_sig00001d9b,
      A3 => blk00000c46_blk00000c47_sig00001d9b,
      CE => ce,
      CLK => clk,
      D => sig00000c23,
      Q => blk00000c46_blk00000c47_sig00001da1,
      Q15 => NLW_blk00000c46_blk00000c47_blk00000c52_Q15_UNCONNECTED
    );
  blk00000c46_blk00000c47_blk00000c51 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000c46_blk00000c47_sig00001da0,
      Q => sig00000c12
    );
  blk00000c46_blk00000c47_blk00000c50 : SRLC16E
    generic map(
      INIT => X"0000"
    )
    port map (
      A0 => blk00000c46_blk00000c47_sig00001d9b,
      A1 => blk00000c46_blk00000c47_sig00001d9c,
      A2 => blk00000c46_blk00000c47_sig00001d9b,
      A3 => blk00000c46_blk00000c47_sig00001d9b,
      CE => ce,
      CLK => clk,
      D => sig00000c20,
      Q => blk00000c46_blk00000c47_sig00001da0,
      Q15 => NLW_blk00000c46_blk00000c47_blk00000c50_Q15_UNCONNECTED
    );
  blk00000c46_blk00000c47_blk00000c4f : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000c46_blk00000c47_sig00001d9f,
      Q => sig00000c11
    );
  blk00000c46_blk00000c47_blk00000c4e : SRLC16E
    generic map(
      INIT => X"0000"
    )
    port map (
      A0 => blk00000c46_blk00000c47_sig00001d9b,
      A1 => blk00000c46_blk00000c47_sig00001d9c,
      A2 => blk00000c46_blk00000c47_sig00001d9b,
      A3 => blk00000c46_blk00000c47_sig00001d9b,
      CE => ce,
      CLK => clk,
      D => sig00000c1f,
      Q => blk00000c46_blk00000c47_sig00001d9f,
      Q15 => NLW_blk00000c46_blk00000c47_blk00000c4e_Q15_UNCONNECTED
    );
  blk00000c46_blk00000c47_blk00000c4d : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000c46_blk00000c47_sig00001d9e,
      Q => sig00000c10
    );
  blk00000c46_blk00000c47_blk00000c4c : SRLC16E
    generic map(
      INIT => X"0000"
    )
    port map (
      A0 => blk00000c46_blk00000c47_sig00001d9b,
      A1 => blk00000c46_blk00000c47_sig00001d9c,
      A2 => blk00000c46_blk00000c47_sig00001d9b,
      A3 => blk00000c46_blk00000c47_sig00001d9b,
      CE => ce,
      CLK => clk,
      D => sig00000c1e,
      Q => blk00000c46_blk00000c47_sig00001d9e,
      Q15 => NLW_blk00000c46_blk00000c47_blk00000c4c_Q15_UNCONNECTED
    );
  blk00000c46_blk00000c47_blk00000c4b : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000c46_blk00000c47_sig00001d9d,
      Q => sig00000c0f
    );
  blk00000c46_blk00000c47_blk00000c4a : SRLC16E
    generic map(
      INIT => X"0000"
    )
    port map (
      A0 => blk00000c46_blk00000c47_sig00001d9b,
      A1 => blk00000c46_blk00000c47_sig00001d9c,
      A2 => blk00000c46_blk00000c47_sig00001d9b,
      A3 => blk00000c46_blk00000c47_sig00001d9b,
      CE => ce,
      CLK => clk,
      D => sig00000c1d,
      Q => blk00000c46_blk00000c47_sig00001d9d,
      Q15 => NLW_blk00000c46_blk00000c47_blk00000c4a_Q15_UNCONNECTED
    );
  blk00000c46_blk00000c47_blk00000c49 : VCC
    port map (
      P => blk00000c46_blk00000c47_sig00001d9c
    );
  blk00000c46_blk00000c47_blk00000c48 : GND
    port map (
      G => blk00000c46_blk00000c47_sig00001d9b
    );
  blk00000c66_blk00000c67_blk00000c85 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000c66_blk00000c67_sig00001df7,
      Q => sig00000a55
    );
  blk00000c66_blk00000c67_blk00000c84 : SRLC16E
    generic map(
      INIT => X"0000"
    )
    port map (
      A0 => blk00000c66_blk00000c67_sig00001de8,
      A1 => blk00000c66_blk00000c67_sig00001de9,
      A2 => blk00000c66_blk00000c67_sig00001de8,
      A3 => blk00000c66_blk00000c67_sig00001de8,
      CE => ce,
      CLK => clk,
      D => sig00000c0d,
      Q => blk00000c66_blk00000c67_sig00001df7,
      Q15 => NLW_blk00000c66_blk00000c67_blk00000c84_Q15_UNCONNECTED
    );
  blk00000c66_blk00000c67_blk00000c83 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000c66_blk00000c67_sig00001df6,
      Q => sig00000a54
    );
  blk00000c66_blk00000c67_blk00000c82 : SRLC16E
    generic map(
      INIT => X"0000"
    )
    port map (
      A0 => blk00000c66_blk00000c67_sig00001de8,
      A1 => blk00000c66_blk00000c67_sig00001de9,
      A2 => blk00000c66_blk00000c67_sig00001de8,
      A3 => blk00000c66_blk00000c67_sig00001de8,
      CE => ce,
      CLK => clk,
      D => sig00000c0c,
      Q => blk00000c66_blk00000c67_sig00001df6,
      Q15 => NLW_blk00000c66_blk00000c67_blk00000c82_Q15_UNCONNECTED
    );
  blk00000c66_blk00000c67_blk00000c81 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000c66_blk00000c67_sig00001df5,
      Q => sig00000a56
    );
  blk00000c66_blk00000c67_blk00000c80 : SRLC16E
    generic map(
      INIT => X"0000"
    )
    port map (
      A0 => blk00000c66_blk00000c67_sig00001de8,
      A1 => blk00000c66_blk00000c67_sig00001de9,
      A2 => blk00000c66_blk00000c67_sig00001de8,
      A3 => blk00000c66_blk00000c67_sig00001de8,
      CE => ce,
      CLK => clk,
      D => sig00000c0e,
      Q => blk00000c66_blk00000c67_sig00001df5,
      Q15 => NLW_blk00000c66_blk00000c67_blk00000c80_Q15_UNCONNECTED
    );
  blk00000c66_blk00000c67_blk00000c7f : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000c66_blk00000c67_sig00001df4,
      Q => sig00000a53
    );
  blk00000c66_blk00000c67_blk00000c7e : SRLC16E
    generic map(
      INIT => X"0000"
    )
    port map (
      A0 => blk00000c66_blk00000c67_sig00001de8,
      A1 => blk00000c66_blk00000c67_sig00001de9,
      A2 => blk00000c66_blk00000c67_sig00001de8,
      A3 => blk00000c66_blk00000c67_sig00001de8,
      CE => ce,
      CLK => clk,
      D => sig00000c0b,
      Q => blk00000c66_blk00000c67_sig00001df4,
      Q15 => NLW_blk00000c66_blk00000c67_blk00000c7e_Q15_UNCONNECTED
    );
  blk00000c66_blk00000c67_blk00000c7d : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000c66_blk00000c67_sig00001df3,
      Q => sig00000a52
    );
  blk00000c66_blk00000c67_blk00000c7c : SRLC16E
    generic map(
      INIT => X"0000"
    )
    port map (
      A0 => blk00000c66_blk00000c67_sig00001de8,
      A1 => blk00000c66_blk00000c67_sig00001de9,
      A2 => blk00000c66_blk00000c67_sig00001de8,
      A3 => blk00000c66_blk00000c67_sig00001de8,
      CE => ce,
      CLK => clk,
      D => sig00000c0a,
      Q => blk00000c66_blk00000c67_sig00001df3,
      Q15 => NLW_blk00000c66_blk00000c67_blk00000c7c_Q15_UNCONNECTED
    );
  blk00000c66_blk00000c67_blk00000c7b : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000c66_blk00000c67_sig00001df2,
      Q => sig00000a51
    );
  blk00000c66_blk00000c67_blk00000c7a : SRLC16E
    generic map(
      INIT => X"0000"
    )
    port map (
      A0 => blk00000c66_blk00000c67_sig00001de8,
      A1 => blk00000c66_blk00000c67_sig00001de9,
      A2 => blk00000c66_blk00000c67_sig00001de8,
      A3 => blk00000c66_blk00000c67_sig00001de8,
      CE => ce,
      CLK => clk,
      D => sig00000c09,
      Q => blk00000c66_blk00000c67_sig00001df2,
      Q15 => NLW_blk00000c66_blk00000c67_blk00000c7a_Q15_UNCONNECTED
    );
  blk00000c66_blk00000c67_blk00000c79 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000c66_blk00000c67_sig00001df1,
      Q => sig00000a50
    );
  blk00000c66_blk00000c67_blk00000c78 : SRLC16E
    generic map(
      INIT => X"0000"
    )
    port map (
      A0 => blk00000c66_blk00000c67_sig00001de8,
      A1 => blk00000c66_blk00000c67_sig00001de9,
      A2 => blk00000c66_blk00000c67_sig00001de8,
      A3 => blk00000c66_blk00000c67_sig00001de8,
      CE => ce,
      CLK => clk,
      D => sig00000c08,
      Q => blk00000c66_blk00000c67_sig00001df1,
      Q15 => NLW_blk00000c66_blk00000c67_blk00000c78_Q15_UNCONNECTED
    );
  blk00000c66_blk00000c67_blk00000c77 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000c66_blk00000c67_sig00001df0,
      Q => sig00000a4e
    );
  blk00000c66_blk00000c67_blk00000c76 : SRLC16E
    generic map(
      INIT => X"0000"
    )
    port map (
      A0 => blk00000c66_blk00000c67_sig00001de8,
      A1 => blk00000c66_blk00000c67_sig00001de9,
      A2 => blk00000c66_blk00000c67_sig00001de8,
      A3 => blk00000c66_blk00000c67_sig00001de8,
      CE => ce,
      CLK => clk,
      D => sig00000c06,
      Q => blk00000c66_blk00000c67_sig00001df0,
      Q15 => NLW_blk00000c66_blk00000c67_blk00000c76_Q15_UNCONNECTED
    );
  blk00000c66_blk00000c67_blk00000c75 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000c66_blk00000c67_sig00001def,
      Q => sig00000a4d
    );
  blk00000c66_blk00000c67_blk00000c74 : SRLC16E
    generic map(
      INIT => X"0000"
    )
    port map (
      A0 => blk00000c66_blk00000c67_sig00001de8,
      A1 => blk00000c66_blk00000c67_sig00001de9,
      A2 => blk00000c66_blk00000c67_sig00001de8,
      A3 => blk00000c66_blk00000c67_sig00001de8,
      CE => ce,
      CLK => clk,
      D => sig00000c05,
      Q => blk00000c66_blk00000c67_sig00001def,
      Q15 => NLW_blk00000c66_blk00000c67_blk00000c74_Q15_UNCONNECTED
    );
  blk00000c66_blk00000c67_blk00000c73 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000c66_blk00000c67_sig00001dee,
      Q => sig00000a4f
    );
  blk00000c66_blk00000c67_blk00000c72 : SRLC16E
    generic map(
      INIT => X"0000"
    )
    port map (
      A0 => blk00000c66_blk00000c67_sig00001de8,
      A1 => blk00000c66_blk00000c67_sig00001de9,
      A2 => blk00000c66_blk00000c67_sig00001de8,
      A3 => blk00000c66_blk00000c67_sig00001de8,
      CE => ce,
      CLK => clk,
      D => sig00000c07,
      Q => blk00000c66_blk00000c67_sig00001dee,
      Q15 => NLW_blk00000c66_blk00000c67_blk00000c72_Q15_UNCONNECTED
    );
  blk00000c66_blk00000c67_blk00000c71 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000c66_blk00000c67_sig00001ded,
      Q => sig00000a4c
    );
  blk00000c66_blk00000c67_blk00000c70 : SRLC16E
    generic map(
      INIT => X"0000"
    )
    port map (
      A0 => blk00000c66_blk00000c67_sig00001de8,
      A1 => blk00000c66_blk00000c67_sig00001de9,
      A2 => blk00000c66_blk00000c67_sig00001de8,
      A3 => blk00000c66_blk00000c67_sig00001de8,
      CE => ce,
      CLK => clk,
      D => sig00000c04,
      Q => blk00000c66_blk00000c67_sig00001ded,
      Q15 => NLW_blk00000c66_blk00000c67_blk00000c70_Q15_UNCONNECTED
    );
  blk00000c66_blk00000c67_blk00000c6f : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000c66_blk00000c67_sig00001dec,
      Q => sig00000a4b
    );
  blk00000c66_blk00000c67_blk00000c6e : SRLC16E
    generic map(
      INIT => X"0000"
    )
    port map (
      A0 => blk00000c66_blk00000c67_sig00001de8,
      A1 => blk00000c66_blk00000c67_sig00001de9,
      A2 => blk00000c66_blk00000c67_sig00001de8,
      A3 => blk00000c66_blk00000c67_sig00001de8,
      CE => ce,
      CLK => clk,
      D => sig00000c03,
      Q => blk00000c66_blk00000c67_sig00001dec,
      Q15 => NLW_blk00000c66_blk00000c67_blk00000c6e_Q15_UNCONNECTED
    );
  blk00000c66_blk00000c67_blk00000c6d : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000c66_blk00000c67_sig00001deb,
      Q => sig00000a4a
    );
  blk00000c66_blk00000c67_blk00000c6c : SRLC16E
    generic map(
      INIT => X"0000"
    )
    port map (
      A0 => blk00000c66_blk00000c67_sig00001de8,
      A1 => blk00000c66_blk00000c67_sig00001de9,
      A2 => blk00000c66_blk00000c67_sig00001de8,
      A3 => blk00000c66_blk00000c67_sig00001de8,
      CE => ce,
      CLK => clk,
      D => sig00000c02,
      Q => blk00000c66_blk00000c67_sig00001deb,
      Q15 => NLW_blk00000c66_blk00000c67_blk00000c6c_Q15_UNCONNECTED
    );
  blk00000c66_blk00000c67_blk00000c6b : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000c66_blk00000c67_sig00001dea,
      Q => sig00000a49
    );
  blk00000c66_blk00000c67_blk00000c6a : SRLC16E
    generic map(
      INIT => X"0000"
    )
    port map (
      A0 => blk00000c66_blk00000c67_sig00001de8,
      A1 => blk00000c66_blk00000c67_sig00001de9,
      A2 => blk00000c66_blk00000c67_sig00001de8,
      A3 => blk00000c66_blk00000c67_sig00001de8,
      CE => ce,
      CLK => clk,
      D => sig00000c01,
      Q => blk00000c66_blk00000c67_sig00001dea,
      Q15 => NLW_blk00000c66_blk00000c67_blk00000c6a_Q15_UNCONNECTED
    );
  blk00000c66_blk00000c67_blk00000c69 : VCC
    port map (
      P => blk00000c66_blk00000c67_sig00001de9
    );
  blk00000c66_blk00000c67_blk00000c68 : GND
    port map (
      G => blk00000c66_blk00000c67_sig00001de8
    );
  blk00000c86_blk00000c87_blk00000c91 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000c86_blk00000c87_sig00001e11,
      Q => sig00000a38
    );
  blk00000c86_blk00000c87_blk00000c90 : SRLC16E
    generic map(
      INIT => X"0000"
    )
    port map (
      A0 => blk00000c86_blk00000c87_sig00001e0c,
      A1 => blk00000c86_blk00000c87_sig00001e0d,
      A2 => blk00000c86_blk00000c87_sig00001e0d,
      A3 => blk00000c86_blk00000c87_sig00001e0d,
      CE => ce,
      CLK => clk,
      D => sig00000a85,
      Q => blk00000c86_blk00000c87_sig00001e11,
      Q15 => NLW_blk00000c86_blk00000c87_blk00000c90_Q15_UNCONNECTED
    );
  blk00000c86_blk00000c87_blk00000c8f : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000c86_blk00000c87_sig00001e10,
      Q => sig00000a37
    );
  blk00000c86_blk00000c87_blk00000c8e : SRLC16E
    generic map(
      INIT => X"0000"
    )
    port map (
      A0 => blk00000c86_blk00000c87_sig00001e0c,
      A1 => blk00000c86_blk00000c87_sig00001e0d,
      A2 => blk00000c86_blk00000c87_sig00001e0d,
      A3 => blk00000c86_blk00000c87_sig00001e0d,
      CE => ce,
      CLK => clk,
      D => sig00000a84,
      Q => blk00000c86_blk00000c87_sig00001e10,
      Q15 => NLW_blk00000c86_blk00000c87_blk00000c8e_Q15_UNCONNECTED
    );
  blk00000c86_blk00000c87_blk00000c8d : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000c86_blk00000c87_sig00001e0f,
      Q => sig00000a3a
    );
  blk00000c86_blk00000c87_blk00000c8c : SRLC16E
    generic map(
      INIT => X"0000"
    )
    port map (
      A0 => blk00000c86_blk00000c87_sig00001e0c,
      A1 => blk00000c86_blk00000c87_sig00001e0d,
      A2 => blk00000c86_blk00000c87_sig00001e0d,
      A3 => blk00000c86_blk00000c87_sig00001e0d,
      CE => ce,
      CLK => clk,
      D => sig00000a83,
      Q => blk00000c86_blk00000c87_sig00001e0f,
      Q15 => NLW_blk00000c86_blk00000c87_blk00000c8c_Q15_UNCONNECTED
    );
  blk00000c86_blk00000c87_blk00000c8b : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000c86_blk00000c87_sig00001e0e,
      Q => sig00000a39
    );
  blk00000c86_blk00000c87_blk00000c8a : SRLC16E
    generic map(
      INIT => X"0000"
    )
    port map (
      A0 => blk00000c86_blk00000c87_sig00001e0c,
      A1 => blk00000c86_blk00000c87_sig00001e0d,
      A2 => blk00000c86_blk00000c87_sig00001e0d,
      A3 => blk00000c86_blk00000c87_sig00001e0d,
      CE => ce,
      CLK => clk,
      D => sig00000a82,
      Q => blk00000c86_blk00000c87_sig00001e0e,
      Q15 => NLW_blk00000c86_blk00000c87_blk00000c8a_Q15_UNCONNECTED
    );
  blk00000c86_blk00000c87_blk00000c89 : VCC
    port map (
      P => blk00000c86_blk00000c87_sig00001e0d
    );
  blk00000c86_blk00000c87_blk00000c88 : GND
    port map (
      G => blk00000c86_blk00000c87_sig00001e0c
    );
  blk00000c92_blk00000c93_blk00000c96 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000c92_blk00000c93_sig00001e22,
      Q => sig00000c96
    );
  blk00000c92_blk00000c93_blk00000c95 : SRLC16E
    generic map(
      INIT => X"0000"
    )
    port map (
      A0 => blk00000c92_blk00000c93_sig00001e21,
      A1 => blk00000c92_blk00000c93_sig00001e21,
      A2 => blk00000c92_blk00000c93_sig00001e21,
      A3 => blk00000c92_blk00000c93_sig00001e21,
      CE => ce,
      CLK => clk,
      D => sig00000c97,
      Q => blk00000c92_blk00000c93_sig00001e22,
      Q15 => NLW_blk00000c92_blk00000c93_blk00000c95_Q15_UNCONNECTED
    );
  blk00000c92_blk00000c93_blk00000c94 : GND
    port map (
      G => blk00000c92_blk00000c93_sig00001e21
    );
  blk00000c9b_blk00000caa : LUT1
    generic map(
      INIT => X"2"
    )
    port map (
      I0 => sig00000a39,
      O => blk00000c9b_sig00001e38
    );
  blk00000c9b_blk00000ca9 : LUT1
    generic map(
      INIT => X"2"
    )
    port map (
      I0 => sig00000a3a,
      O => blk00000c9b_sig00001e37
    );
  blk00000c9b_blk00000ca8 : LUT2
    generic map(
      INIT => X"6"
    )
    port map (
      I0 => sig00000a39,
      I1 => sig00000a3a,
      O => blk00000c9b_sig00001e33
    );
  blk00000c9b_blk00000ca7 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000c9b_sig00001e2f,
      Q => sig00000c9b
    );
  blk00000c9b_blk00000ca6 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000c9b_sig00001e32,
      Q => sig00000c9c
    );
  blk00000c9b_blk00000ca5 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000c9b_sig00001e31,
      Q => sig00000c9d
    );
  blk00000c9b_blk00000ca4 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000c9b_sig00001e30,
      Q => sig00000c9e
    );
  blk00000c9b_blk00000ca3 : MUXCY
    port map (
      CI => blk00000c9b_sig00001e2e,
      DI => sig000008b6,
      S => blk00000c9b_sig00001e38,
      O => blk00000c9b_sig00001e36
    );
  blk00000c9b_blk00000ca2 : MUXCY
    port map (
      CI => blk00000c9b_sig00001e36,
      DI => sig00000a39,
      S => blk00000c9b_sig00001e33,
      O => blk00000c9b_sig00001e35
    );
  blk00000c9b_blk00000ca1 : MUXCY
    port map (
      CI => blk00000c9b_sig00001e35,
      DI => sig00000a3a,
      S => blk00000c9b_sig00001e37,
      O => blk00000c9b_sig00001e34
    );
  blk00000c9b_blk00000ca0 : XORCY
    port map (
      CI => blk00000c9b_sig00001e36,
      LI => blk00000c9b_sig00001e33,
      O => blk00000c9b_sig00001e32
    );
  blk00000c9b_blk00000c9f : XORCY
    port map (
      CI => blk00000c9b_sig00001e35,
      LI => blk00000c9b_sig00001e37,
      O => blk00000c9b_sig00001e31
    );
  blk00000c9b_blk00000c9e : XORCY
    port map (
      CI => blk00000c9b_sig00001e34,
      LI => blk00000c9b_sig00001e2e,
      O => blk00000c9b_sig00001e30
    );
  blk00000c9b_blk00000c9d : XORCY
    port map (
      CI => blk00000c9b_sig00001e2e,
      LI => blk00000c9b_sig00001e38,
      O => blk00000c9b_sig00001e2f
    );
  blk00000c9b_blk00000c9c : GND
    port map (
      G => blk00000c9b_sig00001e2e
    );
  blk00000cb3_blk00000cd5 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000cb3_sig00001e60,
      Q => sig00000a29
    );
  blk00000cb3_blk00000cd4 : SRLC16E
    generic map(
      INIT => X"0000"
    )
    port map (
      A0 => blk00000cb3_sig00001e5e,
      A1 => blk00000cb3_sig00001e5e,
      A2 => blk00000cb3_sig00001e5e,
      A3 => blk00000cb3_sig00001e5e,
      CE => ce,
      CLK => clk,
      D => sig00000c98,
      Q => blk00000cb3_sig00001e60,
      Q15 => NLW_blk00000cb3_blk00000cd4_Q15_UNCONNECTED
    );
  blk00000cb3_blk00000cd3 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000cb3_sig00001e5f,
      Q => sig00000c95
    );
  blk00000cb3_blk00000cd2 : SRLC16E
    generic map(
      INIT => X"0000"
    )
    port map (
      A0 => blk00000cb3_sig00001e5e,
      A1 => blk00000cb3_sig00001e5e,
      A2 => blk00000cb3_sig00001e5e,
      A3 => blk00000cb3_sig00001e5e,
      CE => ce,
      CLK => clk,
      D => sig00000c93,
      Q => blk00000cb3_sig00001e5f,
      Q15 => NLW_blk00000cb3_blk00000cd2_Q15_UNCONNECTED
    );
  blk00000cb3_blk00000cd1 : GND
    port map (
      G => blk00000cb3_sig00001e5e
    );
  blk00000cb3_blk00000cd0 : LUT3
    generic map(
      INIT => X"D8"
    )
    port map (
      I0 => blk00000cb3_sig00001e3f,
      I1 => blk00000cb3_sig00001e4b,
      I2 => blk00000cb3_sig00001e3e,
      O => blk00000cb3_sig00001e53
    );
  blk00000cb3_blk00000ccf : LUT2
    generic map(
      INIT => X"4"
    )
    port map (
      I0 => blk00000cb3_sig00001e3f,
      I1 => blk00000cb3_sig00001e3d,
      O => blk00000cb3_sig00001e52
    );
  blk00000cb3_blk00000cce : LUT3
    generic map(
      INIT => X"D8"
    )
    port map (
      I0 => blk00000cb3_sig00001e3f,
      I1 => blk00000cb3_sig00001e4f,
      I2 => blk00000cb3_sig00001e4d,
      O => blk00000cb3_sig00001e55
    );
  blk00000cb3_blk00000ccd : LUT3
    generic map(
      INIT => X"D8"
    )
    port map (
      I0 => blk00000cb3_sig00001e3f,
      I1 => blk00000cb3_sig00001e4d,
      I2 => blk00000cb3_sig00001e4f,
      O => blk00000cb3_sig00001e54
    );
  blk00000cb3_blk00000ccc : LUT3
    generic map(
      INIT => X"D8"
    )
    port map (
      I0 => blk00000cb3_sig00001e3f,
      I1 => blk00000cb3_sig00001e3e,
      I2 => blk00000cb3_sig00001e4b,
      O => blk00000cb3_sig00001e51
    );
  blk00000cb3_blk00000ccb : LUT2
    generic map(
      INIT => X"8"
    )
    port map (
      I0 => blk00000cb3_sig00001e3f,
      I1 => blk00000cb3_sig00001e3d,
      O => blk00000cb3_sig00001e50
    );
  blk00000cb3_blk00000cca : LUT2
    generic map(
      INIT => X"1"
    )
    port map (
      I0 => sig00000c98,
      I1 => sig00000c99,
      O => blk00000cb3_sig00001e5d
    );
  blk00000cb3_blk00000cc9 : LUT2
    generic map(
      INIT => X"6"
    )
    port map (
      I0 => sig00000c98,
      I1 => sig00000c99,
      O => blk00000cb3_sig00001e5c
    );
  blk00000cb3_blk00000cc8 : LUT2
    generic map(
      INIT => X"E"
    )
    port map (
      I0 => sig00000c99,
      I1 => sig00000c98,
      O => blk00000cb3_sig00001e59
    );
  blk00000cb3_blk00000cc7 : LUT2
    generic map(
      INIT => X"4"
    )
    port map (
      I0 => sig00000c99,
      I1 => sig00000c98,
      O => blk00000cb3_sig00001e58
    );
  blk00000cb3_blk00000cc6 : LUT2
    generic map(
      INIT => X"4"
    )
    port map (
      I0 => sig00000c98,
      I1 => sig00000c99,
      O => blk00000cb3_sig00001e57
    );
  blk00000cb3_blk00000cc5 : LUT2
    generic map(
      INIT => X"8"
    )
    port map (
      I0 => sig00000c98,
      I1 => sig00000c99,
      O => blk00000cb3_sig00001e56
    );
  blk00000cb3_blk00000cc4 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000cb3_sig00001e52,
      Q => sig00000a35
    );
  blk00000cb3_blk00000cc3 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000cb3_sig00001e53,
      Q => sig00000a2f
    );
  blk00000cb3_blk00000cc2 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000cb3_sig00001e50,
      Q => sig00000a2b
    );
  blk00000cb3_blk00000cc1 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000cb3_sig00001e4c,
      Q => sig00000a28
    );
  blk00000cb3_blk00000cc0 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000cb3_sig00001e51,
      Q => sig00000a25
    );
  blk00000cb3_blk00000cbf : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000cb3_sig00001e55,
      Q => sig00000a24
    );
  blk00000cb3_blk00000cbe : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000cb3_sig00001e4e,
      Q => sig00000a23
    );
  blk00000cb3_blk00000cbd : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000cb3_sig00001e54,
      Q => sig00000a22
    );
  blk00000cb3_blk00000cbc : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => sig00000c99,
      Q => blk00000cb3_sig00001e4b
    );
  blk00000cb3_blk00000cbb : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000cb3_sig00001e3f,
      Q => sig00000c94
    );
  blk00000cb3_blk00000cba : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000cb3_sig00001e5d,
      Q => blk00000cb3_sig00001e3d
    );
  blk00000cb3_blk00000cb9 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000cb3_sig00001e59,
      Q => blk00000cb3_sig00001e4c
    );
  blk00000cb3_blk00000cb8 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000cb3_sig00001e5c,
      Q => blk00000cb3_sig00001e3e
    );
  blk00000cb3_blk00000cb7 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000cb3_sig00001e56,
      Q => blk00000cb3_sig00001e4f
    );
  blk00000cb3_blk00000cb6 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000cb3_sig00001e57,
      Q => blk00000cb3_sig00001e4e
    );
  blk00000cb3_blk00000cb5 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000cb3_sig00001e58,
      Q => blk00000cb3_sig00001e4d
    );
  blk00000cb3_blk00000cb4 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => sig00000c9a,
      Q => blk00000cb3_sig00001e3f
    );
  blk00000cd6_blk00000cd7_blk00000ce5 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000cd6_blk00000cd7_sig00001e85,
      Q => sig00000ccf
    );
  blk00000cd6_blk00000cd7_blk00000ce4 : SRLC16E
    generic map(
      INIT => X"0000"
    )
    port map (
      A0 => blk00000cd6_blk00000cd7_sig00001e7f,
      A1 => blk00000cd6_blk00000cd7_sig00001e7e,
      A2 => blk00000cd6_blk00000cd7_sig00001e7e,
      A3 => blk00000cd6_blk00000cd7_sig00001e7e,
      CE => ce,
      CLK => clk,
      D => sig000000e7,
      Q => blk00000cd6_blk00000cd7_sig00001e85,
      Q15 => NLW_blk00000cd6_blk00000cd7_blk00000ce4_Q15_UNCONNECTED
    );
  blk00000cd6_blk00000cd7_blk00000ce3 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000cd6_blk00000cd7_sig00001e84,
      Q => sig00000cce
    );
  blk00000cd6_blk00000cd7_blk00000ce2 : SRLC16E
    generic map(
      INIT => X"0000"
    )
    port map (
      A0 => blk00000cd6_blk00000cd7_sig00001e7f,
      A1 => blk00000cd6_blk00000cd7_sig00001e7e,
      A2 => blk00000cd6_blk00000cd7_sig00001e7e,
      A3 => blk00000cd6_blk00000cd7_sig00001e7e,
      CE => ce,
      CLK => clk,
      D => sig000000e6,
      Q => blk00000cd6_blk00000cd7_sig00001e84,
      Q15 => NLW_blk00000cd6_blk00000cd7_blk00000ce2_Q15_UNCONNECTED
    );
  blk00000cd6_blk00000cd7_blk00000ce1 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000cd6_blk00000cd7_sig00001e83,
      Q => sig00000cd0
    );
  blk00000cd6_blk00000cd7_blk00000ce0 : SRLC16E
    generic map(
      INIT => X"0000"
    )
    port map (
      A0 => blk00000cd6_blk00000cd7_sig00001e7f,
      A1 => blk00000cd6_blk00000cd7_sig00001e7e,
      A2 => blk00000cd6_blk00000cd7_sig00001e7e,
      A3 => blk00000cd6_blk00000cd7_sig00001e7e,
      CE => ce,
      CLK => clk,
      D => sig000000e8,
      Q => blk00000cd6_blk00000cd7_sig00001e83,
      Q15 => NLW_blk00000cd6_blk00000cd7_blk00000ce0_Q15_UNCONNECTED
    );
  blk00000cd6_blk00000cd7_blk00000cdf : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000cd6_blk00000cd7_sig00001e82,
      Q => sig00000ccc
    );
  blk00000cd6_blk00000cd7_blk00000cde : SRLC16E
    generic map(
      INIT => X"0000"
    )
    port map (
      A0 => blk00000cd6_blk00000cd7_sig00001e7f,
      A1 => blk00000cd6_blk00000cd7_sig00001e7e,
      A2 => blk00000cd6_blk00000cd7_sig00001e7e,
      A3 => blk00000cd6_blk00000cd7_sig00001e7e,
      CE => ce,
      CLK => clk,
      D => sig000000e4,
      Q => blk00000cd6_blk00000cd7_sig00001e82,
      Q15 => NLW_blk00000cd6_blk00000cd7_blk00000cde_Q15_UNCONNECTED
    );
  blk00000cd6_blk00000cd7_blk00000cdd : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000cd6_blk00000cd7_sig00001e81,
      Q => sig00000ccb
    );
  blk00000cd6_blk00000cd7_blk00000cdc : SRLC16E
    generic map(
      INIT => X"0000"
    )
    port map (
      A0 => blk00000cd6_blk00000cd7_sig00001e7f,
      A1 => blk00000cd6_blk00000cd7_sig00001e7e,
      A2 => blk00000cd6_blk00000cd7_sig00001e7e,
      A3 => blk00000cd6_blk00000cd7_sig00001e7e,
      CE => ce,
      CLK => clk,
      D => sig000000e3,
      Q => blk00000cd6_blk00000cd7_sig00001e81,
      Q15 => NLW_blk00000cd6_blk00000cd7_blk00000cdc_Q15_UNCONNECTED
    );
  blk00000cd6_blk00000cd7_blk00000cdb : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000cd6_blk00000cd7_sig00001e80,
      Q => sig00000ccd
    );
  blk00000cd6_blk00000cd7_blk00000cda : SRLC16E
    generic map(
      INIT => X"0000"
    )
    port map (
      A0 => blk00000cd6_blk00000cd7_sig00001e7f,
      A1 => blk00000cd6_blk00000cd7_sig00001e7e,
      A2 => blk00000cd6_blk00000cd7_sig00001e7e,
      A3 => blk00000cd6_blk00000cd7_sig00001e7e,
      CE => ce,
      CLK => clk,
      D => sig000000e5,
      Q => blk00000cd6_blk00000cd7_sig00001e80,
      Q15 => NLW_blk00000cd6_blk00000cd7_blk00000cda_Q15_UNCONNECTED
    );
  blk00000cd6_blk00000cd7_blk00000cd9 : VCC
    port map (
      P => blk00000cd6_blk00000cd7_sig00001e7f
    );
  blk00000cd6_blk00000cd7_blk00000cd8 : GND
    port map (
      G => blk00000cd6_blk00000cd7_sig00001e7e
    );
  blk00000ce6_blk00000ce7_blk00000ceb : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000ce6_blk00000ce7_sig00001e97,
      Q => sig00000cca
    );
  blk00000ce6_blk00000ce7_blk00000cea : SRLC16E
    generic map(
      INIT => X"0000"
    )
    port map (
      A0 => blk00000ce6_blk00000ce7_sig00001e96,
      A1 => blk00000ce6_blk00000ce7_sig00001e95,
      A2 => blk00000ce6_blk00000ce7_sig00001e95,
      A3 => blk00000ce6_blk00000ce7_sig00001e95,
      CE => ce,
      CLK => clk,
      D => sig000000ca,
      Q => blk00000ce6_blk00000ce7_sig00001e97,
      Q15 => NLW_blk00000ce6_blk00000ce7_blk00000cea_Q15_UNCONNECTED
    );
  blk00000ce6_blk00000ce7_blk00000ce9 : VCC
    port map (
      P => blk00000ce6_blk00000ce7_sig00001e96
    );
  blk00000ce6_blk00000ce7_blk00000ce8 : GND
    port map (
      G => blk00000ce6_blk00000ce7_sig00001e95
    );
  blk00000cee_blk00000d22 : LUT2
    generic map(
      INIT => X"9"
    )
    port map (
      I0 => sig00000d60,
      I1 => sig00000d7b,
      O => blk00000cee_sig00001ee5
    );
  blk00000cee_blk00000d21 : LUT2
    generic map(
      INIT => X"9"
    )
    port map (
      I0 => sig00000d5e,
      I1 => sig00000d79,
      O => blk00000cee_sig00001ece
    );
  blk00000cee_blk00000d20 : LUT2
    generic map(
      INIT => X"9"
    )
    port map (
      I0 => sig00000d5d,
      I1 => sig00000d78,
      O => blk00000cee_sig00001ecf
    );
  blk00000cee_blk00000d1f : LUT2
    generic map(
      INIT => X"9"
    )
    port map (
      I0 => sig00000d5c,
      I1 => sig00000d77,
      O => blk00000cee_sig00001ed0
    );
  blk00000cee_blk00000d1e : LUT2
    generic map(
      INIT => X"9"
    )
    port map (
      I0 => sig00000d5b,
      I1 => sig00000d76,
      O => blk00000cee_sig00001ed1
    );
  blk00000cee_blk00000d1d : LUT2
    generic map(
      INIT => X"9"
    )
    port map (
      I0 => sig00000d5a,
      I1 => sig00000d75,
      O => blk00000cee_sig00001ed2
    );
  blk00000cee_blk00000d1c : LUT2
    generic map(
      INIT => X"9"
    )
    port map (
      I0 => sig00000d59,
      I1 => sig00000d74,
      O => blk00000cee_sig00001ed3
    );
  blk00000cee_blk00000d1b : LUT2
    generic map(
      INIT => X"9"
    )
    port map (
      I0 => sig00000d58,
      I1 => sig00000d73,
      O => blk00000cee_sig00001ed4
    );
  blk00000cee_blk00000d1a : LUT2
    generic map(
      INIT => X"9"
    )
    port map (
      I0 => sig00000d57,
      I1 => sig00000d72,
      O => blk00000cee_sig00001ed5
    );
  blk00000cee_blk00000d19 : LUT2
    generic map(
      INIT => X"9"
    )
    port map (
      I0 => sig00000d56,
      I1 => sig00000d71,
      O => blk00000cee_sig00001ed6
    );
  blk00000cee_blk00000d18 : LUT2
    generic map(
      INIT => X"9"
    )
    port map (
      I0 => sig00000d60,
      I1 => sig00000d7b,
      O => blk00000cee_sig00001ecc
    );
  blk00000cee_blk00000d17 : LUT2
    generic map(
      INIT => X"9"
    )
    port map (
      I0 => sig00000d5f,
      I1 => sig00000d7a,
      O => blk00000cee_sig00001ecd
    );
  blk00000cee_blk00000d16 : LUT2
    generic map(
      INIT => X"9"
    )
    port map (
      I0 => sig00000d55,
      I1 => sig00000d70,
      O => blk00000cee_sig00001ed7
    );
  blk00000cee_blk00000d15 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000cee_sig00001ecb,
      Q => sig00000d3b
    );
  blk00000cee_blk00000d14 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000cee_sig00001eca,
      Q => sig00000d3c
    );
  blk00000cee_blk00000d13 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000cee_sig00001ec9,
      Q => sig00000d3d
    );
  blk00000cee_blk00000d12 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000cee_sig00001ec8,
      Q => sig00000d3e
    );
  blk00000cee_blk00000d11 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000cee_sig00001ec7,
      Q => sig00000d3f
    );
  blk00000cee_blk00000d10 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000cee_sig00001ec6,
      Q => sig00000d40
    );
  blk00000cee_blk00000d0f : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000cee_sig00001ec5,
      Q => sig00000d41
    );
  blk00000cee_blk00000d0e : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000cee_sig00001ec4,
      Q => sig00000d42
    );
  blk00000cee_blk00000d0d : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000cee_sig00001ec3,
      Q => sig00000d43
    );
  blk00000cee_blk00000d0c : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000cee_sig00001ec2,
      Q => sig00000d44
    );
  blk00000cee_blk00000d0b : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000cee_sig00001ec1,
      Q => sig00000d45
    );
  blk00000cee_blk00000d0a : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000cee_sig00001ec0,
      Q => sig00000d46
    );
  blk00000cee_blk00000d09 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000cee_sig00001ebf,
      Q => sig00000d47
    );
  blk00000cee_blk00000d08 : MUXCY
    port map (
      CI => blk00000cee_sig00001ee4,
      DI => sig00000d55,
      S => blk00000cee_sig00001ed7,
      O => blk00000cee_sig00001ee3
    );
  blk00000cee_blk00000d07 : MUXCY
    port map (
      CI => blk00000cee_sig00001ee3,
      DI => sig00000d56,
      S => blk00000cee_sig00001ed6,
      O => blk00000cee_sig00001ee2
    );
  blk00000cee_blk00000d06 : MUXCY
    port map (
      CI => blk00000cee_sig00001ee2,
      DI => sig00000d57,
      S => blk00000cee_sig00001ed5,
      O => blk00000cee_sig00001ee1
    );
  blk00000cee_blk00000d05 : MUXCY
    port map (
      CI => blk00000cee_sig00001ee1,
      DI => sig00000d58,
      S => blk00000cee_sig00001ed4,
      O => blk00000cee_sig00001ee0
    );
  blk00000cee_blk00000d04 : MUXCY
    port map (
      CI => blk00000cee_sig00001ee0,
      DI => sig00000d59,
      S => blk00000cee_sig00001ed3,
      O => blk00000cee_sig00001edf
    );
  blk00000cee_blk00000d03 : MUXCY
    port map (
      CI => blk00000cee_sig00001edf,
      DI => sig00000d5a,
      S => blk00000cee_sig00001ed2,
      O => blk00000cee_sig00001ede
    );
  blk00000cee_blk00000d02 : MUXCY
    port map (
      CI => blk00000cee_sig00001ede,
      DI => sig00000d5b,
      S => blk00000cee_sig00001ed1,
      O => blk00000cee_sig00001edd
    );
  blk00000cee_blk00000d01 : MUXCY
    port map (
      CI => blk00000cee_sig00001edd,
      DI => sig00000d5c,
      S => blk00000cee_sig00001ed0,
      O => blk00000cee_sig00001edc
    );
  blk00000cee_blk00000d00 : MUXCY
    port map (
      CI => blk00000cee_sig00001edc,
      DI => sig00000d5d,
      S => blk00000cee_sig00001ecf,
      O => blk00000cee_sig00001edb
    );
  blk00000cee_blk00000cff : MUXCY
    port map (
      CI => blk00000cee_sig00001edb,
      DI => sig00000d5e,
      S => blk00000cee_sig00001ece,
      O => blk00000cee_sig00001eda
    );
  blk00000cee_blk00000cfe : MUXCY
    port map (
      CI => blk00000cee_sig00001eda,
      DI => sig00000d5f,
      S => blk00000cee_sig00001ecd,
      O => blk00000cee_sig00001ed9
    );
  blk00000cee_blk00000cfd : MUXCY
    port map (
      CI => blk00000cee_sig00001ed9,
      DI => sig00000d60,
      S => blk00000cee_sig00001ee5,
      O => blk00000cee_sig00001ed8
    );
  blk00000cee_blk00000cfc : XORCY
    port map (
      CI => blk00000cee_sig00001ee4,
      LI => blk00000cee_sig00001ed7,
      O => blk00000cee_sig00001ecb
    );
  blk00000cee_blk00000cfb : XORCY
    port map (
      CI => blk00000cee_sig00001ee3,
      LI => blk00000cee_sig00001ed6,
      O => blk00000cee_sig00001eca
    );
  blk00000cee_blk00000cfa : XORCY
    port map (
      CI => blk00000cee_sig00001ee2,
      LI => blk00000cee_sig00001ed5,
      O => blk00000cee_sig00001ec9
    );
  blk00000cee_blk00000cf9 : XORCY
    port map (
      CI => blk00000cee_sig00001ee1,
      LI => blk00000cee_sig00001ed4,
      O => blk00000cee_sig00001ec8
    );
  blk00000cee_blk00000cf8 : XORCY
    port map (
      CI => blk00000cee_sig00001ee0,
      LI => blk00000cee_sig00001ed3,
      O => blk00000cee_sig00001ec7
    );
  blk00000cee_blk00000cf7 : XORCY
    port map (
      CI => blk00000cee_sig00001edf,
      LI => blk00000cee_sig00001ed2,
      O => blk00000cee_sig00001ec6
    );
  blk00000cee_blk00000cf6 : XORCY
    port map (
      CI => blk00000cee_sig00001ede,
      LI => blk00000cee_sig00001ed1,
      O => blk00000cee_sig00001ec5
    );
  blk00000cee_blk00000cf5 : XORCY
    port map (
      CI => blk00000cee_sig00001edd,
      LI => blk00000cee_sig00001ed0,
      O => blk00000cee_sig00001ec4
    );
  blk00000cee_blk00000cf4 : XORCY
    port map (
      CI => blk00000cee_sig00001edc,
      LI => blk00000cee_sig00001ecf,
      O => blk00000cee_sig00001ec3
    );
  blk00000cee_blk00000cf3 : XORCY
    port map (
      CI => blk00000cee_sig00001edb,
      LI => blk00000cee_sig00001ece,
      O => blk00000cee_sig00001ec2
    );
  blk00000cee_blk00000cf2 : XORCY
    port map (
      CI => blk00000cee_sig00001eda,
      LI => blk00000cee_sig00001ecd,
      O => blk00000cee_sig00001ec1
    );
  blk00000cee_blk00000cf1 : XORCY
    port map (
      CI => blk00000cee_sig00001ed9,
      LI => blk00000cee_sig00001ee5,
      O => blk00000cee_sig00001ec0
    );
  blk00000cee_blk00000cf0 : XORCY
    port map (
      CI => blk00000cee_sig00001ed8,
      LI => blk00000cee_sig00001ecc,
      O => blk00000cee_sig00001ebf
    );
  blk00000cee_blk00000cef : VCC
    port map (
      P => blk00000cee_sig00001ee4
    );
  blk00000d23_blk00000d57 : LUT2
    generic map(
      INIT => X"6"
    )
    port map (
      I0 => sig00000d60,
      I1 => sig00000d7b,
      O => blk00000d23_sig00001f33
    );
  blk00000d23_blk00000d56 : LUT2
    generic map(
      INIT => X"6"
    )
    port map (
      I0 => sig00000d5e,
      I1 => sig00000d79,
      O => blk00000d23_sig00001f1d
    );
  blk00000d23_blk00000d55 : LUT2
    generic map(
      INIT => X"6"
    )
    port map (
      I0 => sig00000d5d,
      I1 => sig00000d78,
      O => blk00000d23_sig00001f1e
    );
  blk00000d23_blk00000d54 : LUT2
    generic map(
      INIT => X"6"
    )
    port map (
      I0 => sig00000d5c,
      I1 => sig00000d77,
      O => blk00000d23_sig00001f1f
    );
  blk00000d23_blk00000d53 : LUT2
    generic map(
      INIT => X"6"
    )
    port map (
      I0 => sig00000d5b,
      I1 => sig00000d76,
      O => blk00000d23_sig00001f20
    );
  blk00000d23_blk00000d52 : LUT2
    generic map(
      INIT => X"6"
    )
    port map (
      I0 => sig00000d5a,
      I1 => sig00000d75,
      O => blk00000d23_sig00001f21
    );
  blk00000d23_blk00000d51 : LUT2
    generic map(
      INIT => X"6"
    )
    port map (
      I0 => sig00000d59,
      I1 => sig00000d74,
      O => blk00000d23_sig00001f22
    );
  blk00000d23_blk00000d50 : LUT2
    generic map(
      INIT => X"6"
    )
    port map (
      I0 => sig00000d58,
      I1 => sig00000d73,
      O => blk00000d23_sig00001f23
    );
  blk00000d23_blk00000d4f : LUT2
    generic map(
      INIT => X"6"
    )
    port map (
      I0 => sig00000d57,
      I1 => sig00000d72,
      O => blk00000d23_sig00001f24
    );
  blk00000d23_blk00000d4e : LUT2
    generic map(
      INIT => X"6"
    )
    port map (
      I0 => sig00000d56,
      I1 => sig00000d71,
      O => blk00000d23_sig00001f25
    );
  blk00000d23_blk00000d4d : LUT2
    generic map(
      INIT => X"6"
    )
    port map (
      I0 => sig00000d60,
      I1 => sig00000d7b,
      O => blk00000d23_sig00001f1b
    );
  blk00000d23_blk00000d4c : LUT2
    generic map(
      INIT => X"6"
    )
    port map (
      I0 => sig00000d5f,
      I1 => sig00000d7a,
      O => blk00000d23_sig00001f1c
    );
  blk00000d23_blk00000d4b : LUT2
    generic map(
      INIT => X"6"
    )
    port map (
      I0 => sig00000d55,
      I1 => sig00000d70,
      O => blk00000d23_sig00001f26
    );
  blk00000d23_blk00000d4a : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000d23_sig00001f1a,
      Q => sig00000d48
    );
  blk00000d23_blk00000d49 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000d23_sig00001f19,
      Q => sig00000d49
    );
  blk00000d23_blk00000d48 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000d23_sig00001f18,
      Q => sig00000d4a
    );
  blk00000d23_blk00000d47 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000d23_sig00001f17,
      Q => sig00000d4b
    );
  blk00000d23_blk00000d46 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000d23_sig00001f16,
      Q => sig00000d4c
    );
  blk00000d23_blk00000d45 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000d23_sig00001f15,
      Q => sig00000d4d
    );
  blk00000d23_blk00000d44 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000d23_sig00001f14,
      Q => sig00000d4e
    );
  blk00000d23_blk00000d43 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000d23_sig00001f13,
      Q => sig00000d4f
    );
  blk00000d23_blk00000d42 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000d23_sig00001f12,
      Q => sig00000d50
    );
  blk00000d23_blk00000d41 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000d23_sig00001f11,
      Q => sig00000d51
    );
  blk00000d23_blk00000d40 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000d23_sig00001f10,
      Q => sig00000d52
    );
  blk00000d23_blk00000d3f : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000d23_sig00001f0f,
      Q => sig00000d53
    );
  blk00000d23_blk00000d3e : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000d23_sig00001f0e,
      Q => sig00000d54
    );
  blk00000d23_blk00000d3d : MUXCY
    port map (
      CI => blk00000d23_sig00001f0d,
      DI => sig00000d55,
      S => blk00000d23_sig00001f26,
      O => blk00000d23_sig00001f32
    );
  blk00000d23_blk00000d3c : MUXCY
    port map (
      CI => blk00000d23_sig00001f32,
      DI => sig00000d56,
      S => blk00000d23_sig00001f25,
      O => blk00000d23_sig00001f31
    );
  blk00000d23_blk00000d3b : MUXCY
    port map (
      CI => blk00000d23_sig00001f31,
      DI => sig00000d57,
      S => blk00000d23_sig00001f24,
      O => blk00000d23_sig00001f30
    );
  blk00000d23_blk00000d3a : MUXCY
    port map (
      CI => blk00000d23_sig00001f30,
      DI => sig00000d58,
      S => blk00000d23_sig00001f23,
      O => blk00000d23_sig00001f2f
    );
  blk00000d23_blk00000d39 : MUXCY
    port map (
      CI => blk00000d23_sig00001f2f,
      DI => sig00000d59,
      S => blk00000d23_sig00001f22,
      O => blk00000d23_sig00001f2e
    );
  blk00000d23_blk00000d38 : MUXCY
    port map (
      CI => blk00000d23_sig00001f2e,
      DI => sig00000d5a,
      S => blk00000d23_sig00001f21,
      O => blk00000d23_sig00001f2d
    );
  blk00000d23_blk00000d37 : MUXCY
    port map (
      CI => blk00000d23_sig00001f2d,
      DI => sig00000d5b,
      S => blk00000d23_sig00001f20,
      O => blk00000d23_sig00001f2c
    );
  blk00000d23_blk00000d36 : MUXCY
    port map (
      CI => blk00000d23_sig00001f2c,
      DI => sig00000d5c,
      S => blk00000d23_sig00001f1f,
      O => blk00000d23_sig00001f2b
    );
  blk00000d23_blk00000d35 : MUXCY
    port map (
      CI => blk00000d23_sig00001f2b,
      DI => sig00000d5d,
      S => blk00000d23_sig00001f1e,
      O => blk00000d23_sig00001f2a
    );
  blk00000d23_blk00000d34 : MUXCY
    port map (
      CI => blk00000d23_sig00001f2a,
      DI => sig00000d5e,
      S => blk00000d23_sig00001f1d,
      O => blk00000d23_sig00001f29
    );
  blk00000d23_blk00000d33 : MUXCY
    port map (
      CI => blk00000d23_sig00001f29,
      DI => sig00000d5f,
      S => blk00000d23_sig00001f1c,
      O => blk00000d23_sig00001f28
    );
  blk00000d23_blk00000d32 : MUXCY
    port map (
      CI => blk00000d23_sig00001f28,
      DI => sig00000d60,
      S => blk00000d23_sig00001f33,
      O => blk00000d23_sig00001f27
    );
  blk00000d23_blk00000d31 : XORCY
    port map (
      CI => blk00000d23_sig00001f0d,
      LI => blk00000d23_sig00001f26,
      O => blk00000d23_sig00001f1a
    );
  blk00000d23_blk00000d30 : XORCY
    port map (
      CI => blk00000d23_sig00001f32,
      LI => blk00000d23_sig00001f25,
      O => blk00000d23_sig00001f19
    );
  blk00000d23_blk00000d2f : XORCY
    port map (
      CI => blk00000d23_sig00001f31,
      LI => blk00000d23_sig00001f24,
      O => blk00000d23_sig00001f18
    );
  blk00000d23_blk00000d2e : XORCY
    port map (
      CI => blk00000d23_sig00001f30,
      LI => blk00000d23_sig00001f23,
      O => blk00000d23_sig00001f17
    );
  blk00000d23_blk00000d2d : XORCY
    port map (
      CI => blk00000d23_sig00001f2f,
      LI => blk00000d23_sig00001f22,
      O => blk00000d23_sig00001f16
    );
  blk00000d23_blk00000d2c : XORCY
    port map (
      CI => blk00000d23_sig00001f2e,
      LI => blk00000d23_sig00001f21,
      O => blk00000d23_sig00001f15
    );
  blk00000d23_blk00000d2b : XORCY
    port map (
      CI => blk00000d23_sig00001f2d,
      LI => blk00000d23_sig00001f20,
      O => blk00000d23_sig00001f14
    );
  blk00000d23_blk00000d2a : XORCY
    port map (
      CI => blk00000d23_sig00001f2c,
      LI => blk00000d23_sig00001f1f,
      O => blk00000d23_sig00001f13
    );
  blk00000d23_blk00000d29 : XORCY
    port map (
      CI => blk00000d23_sig00001f2b,
      LI => blk00000d23_sig00001f1e,
      O => blk00000d23_sig00001f12
    );
  blk00000d23_blk00000d28 : XORCY
    port map (
      CI => blk00000d23_sig00001f2a,
      LI => blk00000d23_sig00001f1d,
      O => blk00000d23_sig00001f11
    );
  blk00000d23_blk00000d27 : XORCY
    port map (
      CI => blk00000d23_sig00001f29,
      LI => blk00000d23_sig00001f1c,
      O => blk00000d23_sig00001f10
    );
  blk00000d23_blk00000d26 : XORCY
    port map (
      CI => blk00000d23_sig00001f28,
      LI => blk00000d23_sig00001f33,
      O => blk00000d23_sig00001f0f
    );
  blk00000d23_blk00000d25 : XORCY
    port map (
      CI => blk00000d23_sig00001f27,
      LI => blk00000d23_sig00001f1b,
      O => blk00000d23_sig00001f0e
    );
  blk00000d23_blk00000d24 : GND
    port map (
      G => blk00000d23_sig00001f0d
    );
  blk00000d58_blk00000d59_blk00000d5c : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000d58_blk00000d59_sig00001f44,
      Q => sig00000d61
    );
  blk00000d58_blk00000d59_blk00000d5b : SRLC16E
    generic map(
      INIT => X"0000"
    )
    port map (
      A0 => blk00000d58_blk00000d59_sig00001f43,
      A1 => blk00000d58_blk00000d59_sig00001f43,
      A2 => blk00000d58_blk00000d59_sig00001f43,
      A3 => blk00000d58_blk00000d59_sig00001f43,
      CE => ce,
      CLK => clk,
      D => sig00000d62,
      Q => blk00000d58_blk00000d59_sig00001f44,
      Q15 => NLW_blk00000d58_blk00000d59_blk00000d5b_Q15_UNCONNECTED
    );
  blk00000d58_blk00000d59_blk00000d5a : GND
    port map (
      G => blk00000d58_blk00000d59_sig00001f43
    );
  blk00000d91_blk00000d92_blk00000dab : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000d91_blk00000d92_sig00001f86,
      Q => sig00000d6e
    );
  blk00000d91_blk00000d92_blk00000daa : SRLC16E
    generic map(
      INIT => X"0000"
    )
    port map (
      A0 => blk00000d91_blk00000d92_sig00001f7a,
      A1 => blk00000d91_blk00000d92_sig00001f7a,
      A2 => blk00000d91_blk00000d92_sig00001f7a,
      A3 => blk00000d91_blk00000d92_sig00001f7a,
      CE => ce,
      CLK => clk,
      D => sig000000d5,
      Q => blk00000d91_blk00000d92_sig00001f86,
      Q15 => NLW_blk00000d91_blk00000d92_blk00000daa_Q15_UNCONNECTED
    );
  blk00000d91_blk00000d92_blk00000da9 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000d91_blk00000d92_sig00001f85,
      Q => sig00000d6d
    );
  blk00000d91_blk00000d92_blk00000da8 : SRLC16E
    generic map(
      INIT => X"0000"
    )
    port map (
      A0 => blk00000d91_blk00000d92_sig00001f7a,
      A1 => blk00000d91_blk00000d92_sig00001f7a,
      A2 => blk00000d91_blk00000d92_sig00001f7a,
      A3 => blk00000d91_blk00000d92_sig00001f7a,
      CE => ce,
      CLK => clk,
      D => sig000000d4,
      Q => blk00000d91_blk00000d92_sig00001f85,
      Q15 => NLW_blk00000d91_blk00000d92_blk00000da8_Q15_UNCONNECTED
    );
  blk00000d91_blk00000d92_blk00000da7 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000d91_blk00000d92_sig00001f84,
      Q => sig00000d6f
    );
  blk00000d91_blk00000d92_blk00000da6 : SRLC16E
    generic map(
      INIT => X"0000"
    )
    port map (
      A0 => blk00000d91_blk00000d92_sig00001f7a,
      A1 => blk00000d91_blk00000d92_sig00001f7a,
      A2 => blk00000d91_blk00000d92_sig00001f7a,
      A3 => blk00000d91_blk00000d92_sig00001f7a,
      CE => ce,
      CLK => clk,
      D => sig000000d6,
      Q => blk00000d91_blk00000d92_sig00001f84,
      Q15 => NLW_blk00000d91_blk00000d92_blk00000da6_Q15_UNCONNECTED
    );
  blk00000d91_blk00000d92_blk00000da5 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000d91_blk00000d92_sig00001f83,
      Q => sig00000d6b
    );
  blk00000d91_blk00000d92_blk00000da4 : SRLC16E
    generic map(
      INIT => X"0000"
    )
    port map (
      A0 => blk00000d91_blk00000d92_sig00001f7a,
      A1 => blk00000d91_blk00000d92_sig00001f7a,
      A2 => blk00000d91_blk00000d92_sig00001f7a,
      A3 => blk00000d91_blk00000d92_sig00001f7a,
      CE => ce,
      CLK => clk,
      D => sig000000d2,
      Q => blk00000d91_blk00000d92_sig00001f83,
      Q15 => NLW_blk00000d91_blk00000d92_blk00000da4_Q15_UNCONNECTED
    );
  blk00000d91_blk00000d92_blk00000da3 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000d91_blk00000d92_sig00001f82,
      Q => sig00000d6a
    );
  blk00000d91_blk00000d92_blk00000da2 : SRLC16E
    generic map(
      INIT => X"0000"
    )
    port map (
      A0 => blk00000d91_blk00000d92_sig00001f7a,
      A1 => blk00000d91_blk00000d92_sig00001f7a,
      A2 => blk00000d91_blk00000d92_sig00001f7a,
      A3 => blk00000d91_blk00000d92_sig00001f7a,
      CE => ce,
      CLK => clk,
      D => sig000000d1,
      Q => blk00000d91_blk00000d92_sig00001f82,
      Q15 => NLW_blk00000d91_blk00000d92_blk00000da2_Q15_UNCONNECTED
    );
  blk00000d91_blk00000d92_blk00000da1 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000d91_blk00000d92_sig00001f81,
      Q => sig00000d6c
    );
  blk00000d91_blk00000d92_blk00000da0 : SRLC16E
    generic map(
      INIT => X"0000"
    )
    port map (
      A0 => blk00000d91_blk00000d92_sig00001f7a,
      A1 => blk00000d91_blk00000d92_sig00001f7a,
      A2 => blk00000d91_blk00000d92_sig00001f7a,
      A3 => blk00000d91_blk00000d92_sig00001f7a,
      CE => ce,
      CLK => clk,
      D => sig000000d3,
      Q => blk00000d91_blk00000d92_sig00001f81,
      Q15 => NLW_blk00000d91_blk00000d92_blk00000da0_Q15_UNCONNECTED
    );
  blk00000d91_blk00000d92_blk00000d9f : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000d91_blk00000d92_sig00001f80,
      Q => sig00000d68
    );
  blk00000d91_blk00000d92_blk00000d9e : SRLC16E
    generic map(
      INIT => X"0000"
    )
    port map (
      A0 => blk00000d91_blk00000d92_sig00001f7a,
      A1 => blk00000d91_blk00000d92_sig00001f7a,
      A2 => blk00000d91_blk00000d92_sig00001f7a,
      A3 => blk00000d91_blk00000d92_sig00001f7a,
      CE => ce,
      CLK => clk,
      D => sig000000cf,
      Q => blk00000d91_blk00000d92_sig00001f80,
      Q15 => NLW_blk00000d91_blk00000d92_blk00000d9e_Q15_UNCONNECTED
    );
  blk00000d91_blk00000d92_blk00000d9d : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000d91_blk00000d92_sig00001f7f,
      Q => sig00000d67
    );
  blk00000d91_blk00000d92_blk00000d9c : SRLC16E
    generic map(
      INIT => X"0000"
    )
    port map (
      A0 => blk00000d91_blk00000d92_sig00001f7a,
      A1 => blk00000d91_blk00000d92_sig00001f7a,
      A2 => blk00000d91_blk00000d92_sig00001f7a,
      A3 => blk00000d91_blk00000d92_sig00001f7a,
      CE => ce,
      CLK => clk,
      D => sig000000ce,
      Q => blk00000d91_blk00000d92_sig00001f7f,
      Q15 => NLW_blk00000d91_blk00000d92_blk00000d9c_Q15_UNCONNECTED
    );
  blk00000d91_blk00000d92_blk00000d9b : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000d91_blk00000d92_sig00001f7e,
      Q => sig00000d69
    );
  blk00000d91_blk00000d92_blk00000d9a : SRLC16E
    generic map(
      INIT => X"0000"
    )
    port map (
      A0 => blk00000d91_blk00000d92_sig00001f7a,
      A1 => blk00000d91_blk00000d92_sig00001f7a,
      A2 => blk00000d91_blk00000d92_sig00001f7a,
      A3 => blk00000d91_blk00000d92_sig00001f7a,
      CE => ce,
      CLK => clk,
      D => sig000000d0,
      Q => blk00000d91_blk00000d92_sig00001f7e,
      Q15 => NLW_blk00000d91_blk00000d92_blk00000d9a_Q15_UNCONNECTED
    );
  blk00000d91_blk00000d92_blk00000d99 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000d91_blk00000d92_sig00001f7d,
      Q => sig00000d65
    );
  blk00000d91_blk00000d92_blk00000d98 : SRLC16E
    generic map(
      INIT => X"0000"
    )
    port map (
      A0 => blk00000d91_blk00000d92_sig00001f7a,
      A1 => blk00000d91_blk00000d92_sig00001f7a,
      A2 => blk00000d91_blk00000d92_sig00001f7a,
      A3 => blk00000d91_blk00000d92_sig00001f7a,
      CE => ce,
      CLK => clk,
      D => sig000000cc,
      Q => blk00000d91_blk00000d92_sig00001f7d,
      Q15 => NLW_blk00000d91_blk00000d92_blk00000d98_Q15_UNCONNECTED
    );
  blk00000d91_blk00000d92_blk00000d97 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000d91_blk00000d92_sig00001f7c,
      Q => sig00000d64
    );
  blk00000d91_blk00000d92_blk00000d96 : SRLC16E
    generic map(
      INIT => X"0000"
    )
    port map (
      A0 => blk00000d91_blk00000d92_sig00001f7a,
      A1 => blk00000d91_blk00000d92_sig00001f7a,
      A2 => blk00000d91_blk00000d92_sig00001f7a,
      A3 => blk00000d91_blk00000d92_sig00001f7a,
      CE => ce,
      CLK => clk,
      D => sig000000cb,
      Q => blk00000d91_blk00000d92_sig00001f7c,
      Q15 => NLW_blk00000d91_blk00000d92_blk00000d96_Q15_UNCONNECTED
    );
  blk00000d91_blk00000d92_blk00000d95 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000d91_blk00000d92_sig00001f7b,
      Q => sig00000d66
    );
  blk00000d91_blk00000d92_blk00000d94 : SRLC16E
    generic map(
      INIT => X"0000"
    )
    port map (
      A0 => blk00000d91_blk00000d92_sig00001f7a,
      A1 => blk00000d91_blk00000d92_sig00001f7a,
      A2 => blk00000d91_blk00000d92_sig00001f7a,
      A3 => blk00000d91_blk00000d92_sig00001f7a,
      CE => ce,
      CLK => clk,
      D => sig000000cd,
      Q => blk00000d91_blk00000d92_sig00001f7b,
      Q15 => NLW_blk00000d91_blk00000d92_blk00000d94_Q15_UNCONNECTED
    );
  blk00000d91_blk00000d92_blk00000d93 : GND
    port map (
      G => blk00000d91_blk00000d92_sig00001f7a
    );
  blk00000dac_blk00000dad_blk00000dc6 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000dac_blk00000dad_sig00001fc8,
      Q => sig00000d5f
    );
  blk00000dac_blk00000dad_blk00000dc5 : SRLC16E
    generic map(
      INIT => X"0000"
    )
    port map (
      A0 => blk00000dac_blk00000dad_sig00001fbc,
      A1 => blk00000dac_blk00000dad_sig00001fbc,
      A2 => blk00000dac_blk00000dad_sig00001fbc,
      A3 => blk00000dac_blk00000dad_sig00001fbc,
      CE => ce,
      CLK => clk,
      D => sig00000d86,
      Q => blk00000dac_blk00000dad_sig00001fc8,
      Q15 => NLW_blk00000dac_blk00000dad_blk00000dc5_Q15_UNCONNECTED
    );
  blk00000dac_blk00000dad_blk00000dc4 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000dac_blk00000dad_sig00001fc7,
      Q => sig00000d5e
    );
  blk00000dac_blk00000dad_blk00000dc3 : SRLC16E
    generic map(
      INIT => X"0000"
    )
    port map (
      A0 => blk00000dac_blk00000dad_sig00001fbc,
      A1 => blk00000dac_blk00000dad_sig00001fbc,
      A2 => blk00000dac_blk00000dad_sig00001fbc,
      A3 => blk00000dac_blk00000dad_sig00001fbc,
      CE => ce,
      CLK => clk,
      D => sig00000d85,
      Q => blk00000dac_blk00000dad_sig00001fc7,
      Q15 => NLW_blk00000dac_blk00000dad_blk00000dc3_Q15_UNCONNECTED
    );
  blk00000dac_blk00000dad_blk00000dc2 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000dac_blk00000dad_sig00001fc6,
      Q => sig00000d60
    );
  blk00000dac_blk00000dad_blk00000dc1 : SRLC16E
    generic map(
      INIT => X"0000"
    )
    port map (
      A0 => blk00000dac_blk00000dad_sig00001fbc,
      A1 => blk00000dac_blk00000dad_sig00001fbc,
      A2 => blk00000dac_blk00000dad_sig00001fbc,
      A3 => blk00000dac_blk00000dad_sig00001fbc,
      CE => ce,
      CLK => clk,
      D => sig00000d87,
      Q => blk00000dac_blk00000dad_sig00001fc6,
      Q15 => NLW_blk00000dac_blk00000dad_blk00000dc1_Q15_UNCONNECTED
    );
  blk00000dac_blk00000dad_blk00000dc0 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000dac_blk00000dad_sig00001fc5,
      Q => sig00000d5c
    );
  blk00000dac_blk00000dad_blk00000dbf : SRLC16E
    generic map(
      INIT => X"0000"
    )
    port map (
      A0 => blk00000dac_blk00000dad_sig00001fbc,
      A1 => blk00000dac_blk00000dad_sig00001fbc,
      A2 => blk00000dac_blk00000dad_sig00001fbc,
      A3 => blk00000dac_blk00000dad_sig00001fbc,
      CE => ce,
      CLK => clk,
      D => sig00000d83,
      Q => blk00000dac_blk00000dad_sig00001fc5,
      Q15 => NLW_blk00000dac_blk00000dad_blk00000dbf_Q15_UNCONNECTED
    );
  blk00000dac_blk00000dad_blk00000dbe : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000dac_blk00000dad_sig00001fc4,
      Q => sig00000d5b
    );
  blk00000dac_blk00000dad_blk00000dbd : SRLC16E
    generic map(
      INIT => X"0000"
    )
    port map (
      A0 => blk00000dac_blk00000dad_sig00001fbc,
      A1 => blk00000dac_blk00000dad_sig00001fbc,
      A2 => blk00000dac_blk00000dad_sig00001fbc,
      A3 => blk00000dac_blk00000dad_sig00001fbc,
      CE => ce,
      CLK => clk,
      D => sig00000d82,
      Q => blk00000dac_blk00000dad_sig00001fc4,
      Q15 => NLW_blk00000dac_blk00000dad_blk00000dbd_Q15_UNCONNECTED
    );
  blk00000dac_blk00000dad_blk00000dbc : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000dac_blk00000dad_sig00001fc3,
      Q => sig00000d5d
    );
  blk00000dac_blk00000dad_blk00000dbb : SRLC16E
    generic map(
      INIT => X"0000"
    )
    port map (
      A0 => blk00000dac_blk00000dad_sig00001fbc,
      A1 => blk00000dac_blk00000dad_sig00001fbc,
      A2 => blk00000dac_blk00000dad_sig00001fbc,
      A3 => blk00000dac_blk00000dad_sig00001fbc,
      CE => ce,
      CLK => clk,
      D => sig00000d84,
      Q => blk00000dac_blk00000dad_sig00001fc3,
      Q15 => NLW_blk00000dac_blk00000dad_blk00000dbb_Q15_UNCONNECTED
    );
  blk00000dac_blk00000dad_blk00000dba : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000dac_blk00000dad_sig00001fc2,
      Q => sig00000d59
    );
  blk00000dac_blk00000dad_blk00000db9 : SRLC16E
    generic map(
      INIT => X"0000"
    )
    port map (
      A0 => blk00000dac_blk00000dad_sig00001fbc,
      A1 => blk00000dac_blk00000dad_sig00001fbc,
      A2 => blk00000dac_blk00000dad_sig00001fbc,
      A3 => blk00000dac_blk00000dad_sig00001fbc,
      CE => ce,
      CLK => clk,
      D => sig00000d80,
      Q => blk00000dac_blk00000dad_sig00001fc2,
      Q15 => NLW_blk00000dac_blk00000dad_blk00000db9_Q15_UNCONNECTED
    );
  blk00000dac_blk00000dad_blk00000db8 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000dac_blk00000dad_sig00001fc1,
      Q => sig00000d58
    );
  blk00000dac_blk00000dad_blk00000db7 : SRLC16E
    generic map(
      INIT => X"0000"
    )
    port map (
      A0 => blk00000dac_blk00000dad_sig00001fbc,
      A1 => blk00000dac_blk00000dad_sig00001fbc,
      A2 => blk00000dac_blk00000dad_sig00001fbc,
      A3 => blk00000dac_blk00000dad_sig00001fbc,
      CE => ce,
      CLK => clk,
      D => sig00000d7f,
      Q => blk00000dac_blk00000dad_sig00001fc1,
      Q15 => NLW_blk00000dac_blk00000dad_blk00000db7_Q15_UNCONNECTED
    );
  blk00000dac_blk00000dad_blk00000db6 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000dac_blk00000dad_sig00001fc0,
      Q => sig00000d5a
    );
  blk00000dac_blk00000dad_blk00000db5 : SRLC16E
    generic map(
      INIT => X"0000"
    )
    port map (
      A0 => blk00000dac_blk00000dad_sig00001fbc,
      A1 => blk00000dac_blk00000dad_sig00001fbc,
      A2 => blk00000dac_blk00000dad_sig00001fbc,
      A3 => blk00000dac_blk00000dad_sig00001fbc,
      CE => ce,
      CLK => clk,
      D => sig00000d81,
      Q => blk00000dac_blk00000dad_sig00001fc0,
      Q15 => NLW_blk00000dac_blk00000dad_blk00000db5_Q15_UNCONNECTED
    );
  blk00000dac_blk00000dad_blk00000db4 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000dac_blk00000dad_sig00001fbf,
      Q => sig00000d56
    );
  blk00000dac_blk00000dad_blk00000db3 : SRLC16E
    generic map(
      INIT => X"0000"
    )
    port map (
      A0 => blk00000dac_blk00000dad_sig00001fbc,
      A1 => blk00000dac_blk00000dad_sig00001fbc,
      A2 => blk00000dac_blk00000dad_sig00001fbc,
      A3 => blk00000dac_blk00000dad_sig00001fbc,
      CE => ce,
      CLK => clk,
      D => sig00000d7d,
      Q => blk00000dac_blk00000dad_sig00001fbf,
      Q15 => NLW_blk00000dac_blk00000dad_blk00000db3_Q15_UNCONNECTED
    );
  blk00000dac_blk00000dad_blk00000db2 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000dac_blk00000dad_sig00001fbe,
      Q => sig00000d55
    );
  blk00000dac_blk00000dad_blk00000db1 : SRLC16E
    generic map(
      INIT => X"0000"
    )
    port map (
      A0 => blk00000dac_blk00000dad_sig00001fbc,
      A1 => blk00000dac_blk00000dad_sig00001fbc,
      A2 => blk00000dac_blk00000dad_sig00001fbc,
      A3 => blk00000dac_blk00000dad_sig00001fbc,
      CE => ce,
      CLK => clk,
      D => sig00000d7c,
      Q => blk00000dac_blk00000dad_sig00001fbe,
      Q15 => NLW_blk00000dac_blk00000dad_blk00000db1_Q15_UNCONNECTED
    );
  blk00000dac_blk00000dad_blk00000db0 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000dac_blk00000dad_sig00001fbd,
      Q => sig00000d57
    );
  blk00000dac_blk00000dad_blk00000daf : SRLC16E
    generic map(
      INIT => X"0000"
    )
    port map (
      A0 => blk00000dac_blk00000dad_sig00001fbc,
      A1 => blk00000dac_blk00000dad_sig00001fbc,
      A2 => blk00000dac_blk00000dad_sig00001fbc,
      A3 => blk00000dac_blk00000dad_sig00001fbc,
      CE => ce,
      CLK => clk,
      D => sig00000d7e,
      Q => blk00000dac_blk00000dad_sig00001fbd,
      Q15 => NLW_blk00000dac_blk00000dad_blk00000daf_Q15_UNCONNECTED
    );
  blk00000dac_blk00000dad_blk00000dae : GND
    port map (
      G => blk00000dac_blk00000dad_sig00001fbc
    );
  blk00000dc7_blk00000dc8_blk00000de3 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000dc7_blk00000dc8_sig0000200f,
      Q => sig00000d39
    );
  blk00000dc7_blk00000dc8_blk00000de2 : SRLC16E
    generic map(
      INIT => X"0000"
    )
    port map (
      A0 => blk00000dc7_blk00000dc8_sig00002002,
      A1 => blk00000dc7_blk00000dc8_sig00002002,
      A2 => blk00000dc7_blk00000dc8_sig00002002,
      A3 => blk00000dc7_blk00000dc8_sig00002002,
      CE => ce,
      CLK => clk,
      D => sig00000d46,
      Q => blk00000dc7_blk00000dc8_sig0000200f,
      Q15 => NLW_blk00000dc7_blk00000dc8_blk00000de2_Q15_UNCONNECTED
    );
  blk00000dc7_blk00000dc8_blk00000de1 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000dc7_blk00000dc8_sig0000200e,
      Q => sig00000d38
    );
  blk00000dc7_blk00000dc8_blk00000de0 : SRLC16E
    generic map(
      INIT => X"0000"
    )
    port map (
      A0 => blk00000dc7_blk00000dc8_sig00002002,
      A1 => blk00000dc7_blk00000dc8_sig00002002,
      A2 => blk00000dc7_blk00000dc8_sig00002002,
      A3 => blk00000dc7_blk00000dc8_sig00002002,
      CE => ce,
      CLK => clk,
      D => sig00000d45,
      Q => blk00000dc7_blk00000dc8_sig0000200e,
      Q15 => NLW_blk00000dc7_blk00000dc8_blk00000de0_Q15_UNCONNECTED
    );
  blk00000dc7_blk00000dc8_blk00000ddf : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000dc7_blk00000dc8_sig0000200d,
      Q => sig00000d3a
    );
  blk00000dc7_blk00000dc8_blk00000dde : SRLC16E
    generic map(
      INIT => X"0000"
    )
    port map (
      A0 => blk00000dc7_blk00000dc8_sig00002002,
      A1 => blk00000dc7_blk00000dc8_sig00002002,
      A2 => blk00000dc7_blk00000dc8_sig00002002,
      A3 => blk00000dc7_blk00000dc8_sig00002002,
      CE => ce,
      CLK => clk,
      D => sig00000d47,
      Q => blk00000dc7_blk00000dc8_sig0000200d,
      Q15 => NLW_blk00000dc7_blk00000dc8_blk00000dde_Q15_UNCONNECTED
    );
  blk00000dc7_blk00000dc8_blk00000ddd : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000dc7_blk00000dc8_sig0000200c,
      Q => sig00000d36
    );
  blk00000dc7_blk00000dc8_blk00000ddc : SRLC16E
    generic map(
      INIT => X"0000"
    )
    port map (
      A0 => blk00000dc7_blk00000dc8_sig00002002,
      A1 => blk00000dc7_blk00000dc8_sig00002002,
      A2 => blk00000dc7_blk00000dc8_sig00002002,
      A3 => blk00000dc7_blk00000dc8_sig00002002,
      CE => ce,
      CLK => clk,
      D => sig00000d43,
      Q => blk00000dc7_blk00000dc8_sig0000200c,
      Q15 => NLW_blk00000dc7_blk00000dc8_blk00000ddc_Q15_UNCONNECTED
    );
  blk00000dc7_blk00000dc8_blk00000ddb : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000dc7_blk00000dc8_sig0000200b,
      Q => sig00000d35
    );
  blk00000dc7_blk00000dc8_blk00000dda : SRLC16E
    generic map(
      INIT => X"0000"
    )
    port map (
      A0 => blk00000dc7_blk00000dc8_sig00002002,
      A1 => blk00000dc7_blk00000dc8_sig00002002,
      A2 => blk00000dc7_blk00000dc8_sig00002002,
      A3 => blk00000dc7_blk00000dc8_sig00002002,
      CE => ce,
      CLK => clk,
      D => sig00000d42,
      Q => blk00000dc7_blk00000dc8_sig0000200b,
      Q15 => NLW_blk00000dc7_blk00000dc8_blk00000dda_Q15_UNCONNECTED
    );
  blk00000dc7_blk00000dc8_blk00000dd9 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000dc7_blk00000dc8_sig0000200a,
      Q => sig00000d37
    );
  blk00000dc7_blk00000dc8_blk00000dd8 : SRLC16E
    generic map(
      INIT => X"0000"
    )
    port map (
      A0 => blk00000dc7_blk00000dc8_sig00002002,
      A1 => blk00000dc7_blk00000dc8_sig00002002,
      A2 => blk00000dc7_blk00000dc8_sig00002002,
      A3 => blk00000dc7_blk00000dc8_sig00002002,
      CE => ce,
      CLK => clk,
      D => sig00000d44,
      Q => blk00000dc7_blk00000dc8_sig0000200a,
      Q15 => NLW_blk00000dc7_blk00000dc8_blk00000dd8_Q15_UNCONNECTED
    );
  blk00000dc7_blk00000dc8_blk00000dd7 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000dc7_blk00000dc8_sig00002009,
      Q => sig00000d33
    );
  blk00000dc7_blk00000dc8_blk00000dd6 : SRLC16E
    generic map(
      INIT => X"0000"
    )
    port map (
      A0 => blk00000dc7_blk00000dc8_sig00002002,
      A1 => blk00000dc7_blk00000dc8_sig00002002,
      A2 => blk00000dc7_blk00000dc8_sig00002002,
      A3 => blk00000dc7_blk00000dc8_sig00002002,
      CE => ce,
      CLK => clk,
      D => sig00000d40,
      Q => blk00000dc7_blk00000dc8_sig00002009,
      Q15 => NLW_blk00000dc7_blk00000dc8_blk00000dd6_Q15_UNCONNECTED
    );
  blk00000dc7_blk00000dc8_blk00000dd5 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000dc7_blk00000dc8_sig00002008,
      Q => sig00000d32
    );
  blk00000dc7_blk00000dc8_blk00000dd4 : SRLC16E
    generic map(
      INIT => X"0000"
    )
    port map (
      A0 => blk00000dc7_blk00000dc8_sig00002002,
      A1 => blk00000dc7_blk00000dc8_sig00002002,
      A2 => blk00000dc7_blk00000dc8_sig00002002,
      A3 => blk00000dc7_blk00000dc8_sig00002002,
      CE => ce,
      CLK => clk,
      D => sig00000d3f,
      Q => blk00000dc7_blk00000dc8_sig00002008,
      Q15 => NLW_blk00000dc7_blk00000dc8_blk00000dd4_Q15_UNCONNECTED
    );
  blk00000dc7_blk00000dc8_blk00000dd3 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000dc7_blk00000dc8_sig00002007,
      Q => sig00000d34
    );
  blk00000dc7_blk00000dc8_blk00000dd2 : SRLC16E
    generic map(
      INIT => X"0000"
    )
    port map (
      A0 => blk00000dc7_blk00000dc8_sig00002002,
      A1 => blk00000dc7_blk00000dc8_sig00002002,
      A2 => blk00000dc7_blk00000dc8_sig00002002,
      A3 => blk00000dc7_blk00000dc8_sig00002002,
      CE => ce,
      CLK => clk,
      D => sig00000d41,
      Q => blk00000dc7_blk00000dc8_sig00002007,
      Q15 => NLW_blk00000dc7_blk00000dc8_blk00000dd2_Q15_UNCONNECTED
    );
  blk00000dc7_blk00000dc8_blk00000dd1 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000dc7_blk00000dc8_sig00002006,
      Q => sig00000d31
    );
  blk00000dc7_blk00000dc8_blk00000dd0 : SRLC16E
    generic map(
      INIT => X"0000"
    )
    port map (
      A0 => blk00000dc7_blk00000dc8_sig00002002,
      A1 => blk00000dc7_blk00000dc8_sig00002002,
      A2 => blk00000dc7_blk00000dc8_sig00002002,
      A3 => blk00000dc7_blk00000dc8_sig00002002,
      CE => ce,
      CLK => clk,
      D => sig00000d3e,
      Q => blk00000dc7_blk00000dc8_sig00002006,
      Q15 => NLW_blk00000dc7_blk00000dc8_blk00000dd0_Q15_UNCONNECTED
    );
  blk00000dc7_blk00000dc8_blk00000dcf : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000dc7_blk00000dc8_sig00002005,
      Q => sig00000d30
    );
  blk00000dc7_blk00000dc8_blk00000dce : SRLC16E
    generic map(
      INIT => X"0000"
    )
    port map (
      A0 => blk00000dc7_blk00000dc8_sig00002002,
      A1 => blk00000dc7_blk00000dc8_sig00002002,
      A2 => blk00000dc7_blk00000dc8_sig00002002,
      A3 => blk00000dc7_blk00000dc8_sig00002002,
      CE => ce,
      CLK => clk,
      D => sig00000d3d,
      Q => blk00000dc7_blk00000dc8_sig00002005,
      Q15 => NLW_blk00000dc7_blk00000dc8_blk00000dce_Q15_UNCONNECTED
    );
  blk00000dc7_blk00000dc8_blk00000dcd : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000dc7_blk00000dc8_sig00002004,
      Q => sig00000d2f
    );
  blk00000dc7_blk00000dc8_blk00000dcc : SRLC16E
    generic map(
      INIT => X"0000"
    )
    port map (
      A0 => blk00000dc7_blk00000dc8_sig00002002,
      A1 => blk00000dc7_blk00000dc8_sig00002002,
      A2 => blk00000dc7_blk00000dc8_sig00002002,
      A3 => blk00000dc7_blk00000dc8_sig00002002,
      CE => ce,
      CLK => clk,
      D => sig00000d3c,
      Q => blk00000dc7_blk00000dc8_sig00002004,
      Q15 => NLW_blk00000dc7_blk00000dc8_blk00000dcc_Q15_UNCONNECTED
    );
  blk00000dc7_blk00000dc8_blk00000dcb : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000dc7_blk00000dc8_sig00002003,
      Q => sig00000d2e
    );
  blk00000dc7_blk00000dc8_blk00000dca : SRLC16E
    generic map(
      INIT => X"0000"
    )
    port map (
      A0 => blk00000dc7_blk00000dc8_sig00002002,
      A1 => blk00000dc7_blk00000dc8_sig00002002,
      A2 => blk00000dc7_blk00000dc8_sig00002002,
      A3 => blk00000dc7_blk00000dc8_sig00002002,
      CE => ce,
      CLK => clk,
      D => sig00000d3b,
      Q => blk00000dc7_blk00000dc8_sig00002003,
      Q15 => NLW_blk00000dc7_blk00000dc8_blk00000dca_Q15_UNCONNECTED
    );
  blk00000dc7_blk00000dc8_blk00000dc9 : GND
    port map (
      G => blk00000dc7_blk00000dc8_sig00002002
    );
  blk00000de4_blk00000de5_blk00000e00 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000de4_blk00000de5_sig00002056,
      Q => sig00000ced
    );
  blk00000de4_blk00000de5_blk00000dff : SRLC16E
    generic map(
      INIT => X"0000"
    )
    port map (
      A0 => blk00000de4_blk00000de5_sig00002049,
      A1 => blk00000de4_blk00000de5_sig00002049,
      A2 => blk00000de4_blk00000de5_sig00002049,
      A3 => blk00000de4_blk00000de5_sig00002049,
      CE => ce,
      CLK => clk,
      D => sig00000d2c,
      Q => blk00000de4_blk00000de5_sig00002056,
      Q15 => NLW_blk00000de4_blk00000de5_blk00000dff_Q15_UNCONNECTED
    );
  blk00000de4_blk00000de5_blk00000dfe : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000de4_blk00000de5_sig00002055,
      Q => sig00000cec
    );
  blk00000de4_blk00000de5_blk00000dfd : SRLC16E
    generic map(
      INIT => X"0000"
    )
    port map (
      A0 => blk00000de4_blk00000de5_sig00002049,
      A1 => blk00000de4_blk00000de5_sig00002049,
      A2 => blk00000de4_blk00000de5_sig00002049,
      A3 => blk00000de4_blk00000de5_sig00002049,
      CE => ce,
      CLK => clk,
      D => sig00000d2b,
      Q => blk00000de4_blk00000de5_sig00002055,
      Q15 => NLW_blk00000de4_blk00000de5_blk00000dfd_Q15_UNCONNECTED
    );
  blk00000de4_blk00000de5_blk00000dfc : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000de4_blk00000de5_sig00002054,
      Q => sig00000cee
    );
  blk00000de4_blk00000de5_blk00000dfb : SRLC16E
    generic map(
      INIT => X"0000"
    )
    port map (
      A0 => blk00000de4_blk00000de5_sig00002049,
      A1 => blk00000de4_blk00000de5_sig00002049,
      A2 => blk00000de4_blk00000de5_sig00002049,
      A3 => blk00000de4_blk00000de5_sig00002049,
      CE => ce,
      CLK => clk,
      D => sig00000d2d,
      Q => blk00000de4_blk00000de5_sig00002054,
      Q15 => NLW_blk00000de4_blk00000de5_blk00000dfb_Q15_UNCONNECTED
    );
  blk00000de4_blk00000de5_blk00000dfa : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000de4_blk00000de5_sig00002053,
      Q => sig00000cea
    );
  blk00000de4_blk00000de5_blk00000df9 : SRLC16E
    generic map(
      INIT => X"0000"
    )
    port map (
      A0 => blk00000de4_blk00000de5_sig00002049,
      A1 => blk00000de4_blk00000de5_sig00002049,
      A2 => blk00000de4_blk00000de5_sig00002049,
      A3 => blk00000de4_blk00000de5_sig00002049,
      CE => ce,
      CLK => clk,
      D => sig00000d29,
      Q => blk00000de4_blk00000de5_sig00002053,
      Q15 => NLW_blk00000de4_blk00000de5_blk00000df9_Q15_UNCONNECTED
    );
  blk00000de4_blk00000de5_blk00000df8 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000de4_blk00000de5_sig00002052,
      Q => sig00000ce9
    );
  blk00000de4_blk00000de5_blk00000df7 : SRLC16E
    generic map(
      INIT => X"0000"
    )
    port map (
      A0 => blk00000de4_blk00000de5_sig00002049,
      A1 => blk00000de4_blk00000de5_sig00002049,
      A2 => blk00000de4_blk00000de5_sig00002049,
      A3 => blk00000de4_blk00000de5_sig00002049,
      CE => ce,
      CLK => clk,
      D => sig00000d28,
      Q => blk00000de4_blk00000de5_sig00002052,
      Q15 => NLW_blk00000de4_blk00000de5_blk00000df7_Q15_UNCONNECTED
    );
  blk00000de4_blk00000de5_blk00000df6 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000de4_blk00000de5_sig00002051,
      Q => sig00000ceb
    );
  blk00000de4_blk00000de5_blk00000df5 : SRLC16E
    generic map(
      INIT => X"0000"
    )
    port map (
      A0 => blk00000de4_blk00000de5_sig00002049,
      A1 => blk00000de4_blk00000de5_sig00002049,
      A2 => blk00000de4_blk00000de5_sig00002049,
      A3 => blk00000de4_blk00000de5_sig00002049,
      CE => ce,
      CLK => clk,
      D => sig00000d2a,
      Q => blk00000de4_blk00000de5_sig00002051,
      Q15 => NLW_blk00000de4_blk00000de5_blk00000df5_Q15_UNCONNECTED
    );
  blk00000de4_blk00000de5_blk00000df4 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000de4_blk00000de5_sig00002050,
      Q => sig00000ce7
    );
  blk00000de4_blk00000de5_blk00000df3 : SRLC16E
    generic map(
      INIT => X"0000"
    )
    port map (
      A0 => blk00000de4_blk00000de5_sig00002049,
      A1 => blk00000de4_blk00000de5_sig00002049,
      A2 => blk00000de4_blk00000de5_sig00002049,
      A3 => blk00000de4_blk00000de5_sig00002049,
      CE => ce,
      CLK => clk,
      D => sig00000d26,
      Q => blk00000de4_blk00000de5_sig00002050,
      Q15 => NLW_blk00000de4_blk00000de5_blk00000df3_Q15_UNCONNECTED
    );
  blk00000de4_blk00000de5_blk00000df2 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000de4_blk00000de5_sig0000204f,
      Q => sig00000ce6
    );
  blk00000de4_blk00000de5_blk00000df1 : SRLC16E
    generic map(
      INIT => X"0000"
    )
    port map (
      A0 => blk00000de4_blk00000de5_sig00002049,
      A1 => blk00000de4_blk00000de5_sig00002049,
      A2 => blk00000de4_blk00000de5_sig00002049,
      A3 => blk00000de4_blk00000de5_sig00002049,
      CE => ce,
      CLK => clk,
      D => sig00000d25,
      Q => blk00000de4_blk00000de5_sig0000204f,
      Q15 => NLW_blk00000de4_blk00000de5_blk00000df1_Q15_UNCONNECTED
    );
  blk00000de4_blk00000de5_blk00000df0 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000de4_blk00000de5_sig0000204e,
      Q => sig00000ce8
    );
  blk00000de4_blk00000de5_blk00000def : SRLC16E
    generic map(
      INIT => X"0000"
    )
    port map (
      A0 => blk00000de4_blk00000de5_sig00002049,
      A1 => blk00000de4_blk00000de5_sig00002049,
      A2 => blk00000de4_blk00000de5_sig00002049,
      A3 => blk00000de4_blk00000de5_sig00002049,
      CE => ce,
      CLK => clk,
      D => sig00000d27,
      Q => blk00000de4_blk00000de5_sig0000204e,
      Q15 => NLW_blk00000de4_blk00000de5_blk00000def_Q15_UNCONNECTED
    );
  blk00000de4_blk00000de5_blk00000dee : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000de4_blk00000de5_sig0000204d,
      Q => sig00000ce5
    );
  blk00000de4_blk00000de5_blk00000ded : SRLC16E
    generic map(
      INIT => X"0000"
    )
    port map (
      A0 => blk00000de4_blk00000de5_sig00002049,
      A1 => blk00000de4_blk00000de5_sig00002049,
      A2 => blk00000de4_blk00000de5_sig00002049,
      A3 => blk00000de4_blk00000de5_sig00002049,
      CE => ce,
      CLK => clk,
      D => sig00000d24,
      Q => blk00000de4_blk00000de5_sig0000204d,
      Q15 => NLW_blk00000de4_blk00000de5_blk00000ded_Q15_UNCONNECTED
    );
  blk00000de4_blk00000de5_blk00000dec : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000de4_blk00000de5_sig0000204c,
      Q => sig00000ce4
    );
  blk00000de4_blk00000de5_blk00000deb : SRLC16E
    generic map(
      INIT => X"0000"
    )
    port map (
      A0 => blk00000de4_blk00000de5_sig00002049,
      A1 => blk00000de4_blk00000de5_sig00002049,
      A2 => blk00000de4_blk00000de5_sig00002049,
      A3 => blk00000de4_blk00000de5_sig00002049,
      CE => ce,
      CLK => clk,
      D => sig00000d23,
      Q => blk00000de4_blk00000de5_sig0000204c,
      Q15 => NLW_blk00000de4_blk00000de5_blk00000deb_Q15_UNCONNECTED
    );
  blk00000de4_blk00000de5_blk00000dea : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000de4_blk00000de5_sig0000204b,
      Q => sig00000ce3
    );
  blk00000de4_blk00000de5_blk00000de9 : SRLC16E
    generic map(
      INIT => X"0000"
    )
    port map (
      A0 => blk00000de4_blk00000de5_sig00002049,
      A1 => blk00000de4_blk00000de5_sig00002049,
      A2 => blk00000de4_blk00000de5_sig00002049,
      A3 => blk00000de4_blk00000de5_sig00002049,
      CE => ce,
      CLK => clk,
      D => sig00000d22,
      Q => blk00000de4_blk00000de5_sig0000204b,
      Q15 => NLW_blk00000de4_blk00000de5_blk00000de9_Q15_UNCONNECTED
    );
  blk00000de4_blk00000de5_blk00000de8 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000de4_blk00000de5_sig0000204a,
      Q => sig00000ce2
    );
  blk00000de4_blk00000de5_blk00000de7 : SRLC16E
    generic map(
      INIT => X"0000"
    )
    port map (
      A0 => blk00000de4_blk00000de5_sig00002049,
      A1 => blk00000de4_blk00000de5_sig00002049,
      A2 => blk00000de4_blk00000de5_sig00002049,
      A3 => blk00000de4_blk00000de5_sig00002049,
      CE => ce,
      CLK => clk,
      D => sig00000d21,
      Q => blk00000de4_blk00000de5_sig0000204a,
      Q15 => NLW_blk00000de4_blk00000de5_blk00000de7_Q15_UNCONNECTED
    );
  blk00000de4_blk00000de5_blk00000de6 : GND
    port map (
      G => blk00000de4_blk00000de5_sig00002049
    );
  blk00000e01_blk00000e02_blk00000e08 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000e01_blk00000e02_sig00002066,
      Q => sig00000cd4
    );
  blk00000e01_blk00000e02_blk00000e07 : SRLC16E
    generic map(
      INIT => X"0000"
    )
    port map (
      A0 => blk00000e01_blk00000e02_sig00002063,
      A1 => blk00000e01_blk00000e02_sig00002063,
      A2 => blk00000e01_blk00000e02_sig00002064,
      A3 => blk00000e01_blk00000e02_sig00002063,
      CE => ce,
      CLK => clk,
      D => sig000000ec,
      Q => blk00000e01_blk00000e02_sig00002066,
      Q15 => NLW_blk00000e01_blk00000e02_blk00000e07_Q15_UNCONNECTED
    );
  blk00000e01_blk00000e02_blk00000e06 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000e01_blk00000e02_sig00002065,
      Q => sig00000cd3
    );
  blk00000e01_blk00000e02_blk00000e05 : SRLC16E
    generic map(
      INIT => X"0000"
    )
    port map (
      A0 => blk00000e01_blk00000e02_sig00002063,
      A1 => blk00000e01_blk00000e02_sig00002063,
      A2 => blk00000e01_blk00000e02_sig00002064,
      A3 => blk00000e01_blk00000e02_sig00002063,
      CE => ce,
      CLK => clk,
      D => sig000000eb,
      Q => blk00000e01_blk00000e02_sig00002065,
      Q15 => NLW_blk00000e01_blk00000e02_blk00000e05_Q15_UNCONNECTED
    );
  blk00000e01_blk00000e02_blk00000e04 : VCC
    port map (
      P => blk00000e01_blk00000e02_sig00002064
    );
  blk00000e01_blk00000e02_blk00000e03 : GND
    port map (
      G => blk00000e01_blk00000e02_sig00002063
    );
  blk00000e09_blk00000e0a_blk00000e10 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000e09_blk00000e0a_sig00002076,
      Q => sig00000cd2
    );
  blk00000e09_blk00000e0a_blk00000e0f : SRLC16E
    generic map(
      INIT => X"0000"
    )
    port map (
      A0 => blk00000e09_blk00000e0a_sig00002074,
      A1 => blk00000e09_blk00000e0a_sig00002073,
      A2 => blk00000e09_blk00000e0a_sig00002073,
      A3 => blk00000e09_blk00000e0a_sig00002073,
      CE => ce,
      CLK => clk,
      D => sig000000ea,
      Q => blk00000e09_blk00000e0a_sig00002076,
      Q15 => NLW_blk00000e09_blk00000e0a_blk00000e0f_Q15_UNCONNECTED
    );
  blk00000e09_blk00000e0a_blk00000e0e : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000e09_blk00000e0a_sig00002075,
      Q => sig00000cd1
    );
  blk00000e09_blk00000e0a_blk00000e0d : SRLC16E
    generic map(
      INIT => X"0000"
    )
    port map (
      A0 => blk00000e09_blk00000e0a_sig00002074,
      A1 => blk00000e09_blk00000e0a_sig00002073,
      A2 => blk00000e09_blk00000e0a_sig00002073,
      A3 => blk00000e09_blk00000e0a_sig00002073,
      CE => ce,
      CLK => clk,
      D => sig000000e9,
      Q => blk00000e09_blk00000e0a_sig00002075,
      Q15 => NLW_blk00000e09_blk00000e0a_blk00000e0d_Q15_UNCONNECTED
    );
  blk00000e09_blk00000e0a_blk00000e0c : VCC
    port map (
      P => blk00000e09_blk00000e0a_sig00002074
    );
  blk00000e09_blk00000e0a_blk00000e0b : GND
    port map (
      G => blk00000e09_blk00000e0a_sig00002073
    );
  blk00000e11_blk00000e12_blk00000e16 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000e11_blk00000e12_sig00002081,
      Q => sig00000ca7
    );
  blk00000e11_blk00000e12_blk00000e15 : SRLC16E
    generic map(
      INIT => X"0000"
    )
    port map (
      A0 => blk00000e11_blk00000e12_sig00002080,
      A1 => blk00000e11_blk00000e12_sig00002080,
      A2 => blk00000e11_blk00000e12_sig00002080,
      A3 => blk00000e11_blk00000e12_sig0000207f,
      CE => ce,
      CLK => clk,
      D => sig00000cca,
      Q => blk00000e11_blk00000e12_sig00002081,
      Q15 => NLW_blk00000e11_blk00000e12_blk00000e15_Q15_UNCONNECTED
    );
  blk00000e11_blk00000e12_blk00000e14 : VCC
    port map (
      P => blk00000e11_blk00000e12_sig00002080
    );
  blk00000e11_blk00000e12_blk00000e13 : GND
    port map (
      G => blk00000e11_blk00000e12_sig0000207f
    );
  blk00000e17_blk00000e18_blk00000e1c : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000e17_blk00000e18_sig0000208c,
      Q => sig00000cc8
    );
  blk00000e17_blk00000e18_blk00000e1b : SRLC16E
    generic map(
      INIT => X"0000"
    )
    port map (
      A0 => blk00000e17_blk00000e18_sig0000208b,
      A1 => blk00000e17_blk00000e18_sig0000208b,
      A2 => blk00000e17_blk00000e18_sig0000208a,
      A3 => blk00000e17_blk00000e18_sig0000208a,
      CE => ce,
      CLK => clk,
      D => sig00000cc9,
      Q => blk00000e17_blk00000e18_sig0000208c,
      Q15 => NLW_blk00000e17_blk00000e18_blk00000e1b_Q15_UNCONNECTED
    );
  blk00000e17_blk00000e18_blk00000e1a : VCC
    port map (
      P => blk00000e17_blk00000e18_sig0000208b
    );
  blk00000e17_blk00000e18_blk00000e19 : GND
    port map (
      G => blk00000e17_blk00000e18_sig0000208a
    );
  blk00000e1d_blk00000e1e_blk00000e24 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000e1d_blk00000e1e_sig0000209c,
      Q => sig00000cc7
    );
  blk00000e1d_blk00000e1e_blk00000e23 : SRLC16E
    generic map(
      INIT => X"0000"
    )
    port map (
      A0 => blk00000e1d_blk00000e1e_sig0000209a,
      A1 => blk00000e1d_blk00000e1e_sig00002099,
      A2 => blk00000e1d_blk00000e1e_sig00002099,
      A3 => blk00000e1d_blk00000e1e_sig0000209a,
      CE => ce,
      CLK => clk,
      D => sig00000cd2,
      Q => blk00000e1d_blk00000e1e_sig0000209c,
      Q15 => NLW_blk00000e1d_blk00000e1e_blk00000e23_Q15_UNCONNECTED
    );
  blk00000e1d_blk00000e1e_blk00000e22 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000e1d_blk00000e1e_sig0000209b,
      Q => sig00000cc6
    );
  blk00000e1d_blk00000e1e_blk00000e21 : SRLC16E
    generic map(
      INIT => X"0000"
    )
    port map (
      A0 => blk00000e1d_blk00000e1e_sig0000209a,
      A1 => blk00000e1d_blk00000e1e_sig00002099,
      A2 => blk00000e1d_blk00000e1e_sig00002099,
      A3 => blk00000e1d_blk00000e1e_sig0000209a,
      CE => ce,
      CLK => clk,
      D => sig00000cd1,
      Q => blk00000e1d_blk00000e1e_sig0000209b,
      Q15 => NLW_blk00000e1d_blk00000e1e_blk00000e21_Q15_UNCONNECTED
    );
  blk00000e1d_blk00000e1e_blk00000e20 : VCC
    port map (
      P => blk00000e1d_blk00000e1e_sig0000209a
    );
  blk00000e1d_blk00000e1e_blk00000e1f : GND
    port map (
      G => blk00000e1d_blk00000e1e_sig00002099
    );
  blk00000e25_blk00000e26_blk00000e34 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000e25_blk00000e26_sig000020c0,
      Q => sig000000c7
    );
  blk00000e25_blk00000e26_blk00000e33 : SRLC16E
    generic map(
      INIT => X"0000"
    )
    port map (
      A0 => blk00000e25_blk00000e26_sig000020b9,
      A1 => blk00000e25_blk00000e26_sig000020ba,
      A2 => blk00000e25_blk00000e26_sig000020b9,
      A3 => blk00000e25_blk00000e26_sig000020ba,
      CE => ce,
      CLK => clk,
      D => sig00000ccf,
      Q => blk00000e25_blk00000e26_sig000020c0,
      Q15 => NLW_blk00000e25_blk00000e26_blk00000e33_Q15_UNCONNECTED
    );
  blk00000e25_blk00000e26_blk00000e32 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000e25_blk00000e26_sig000020bf,
      Q => sig000000c6
    );
  blk00000e25_blk00000e26_blk00000e31 : SRLC16E
    generic map(
      INIT => X"0000"
    )
    port map (
      A0 => blk00000e25_blk00000e26_sig000020b9,
      A1 => blk00000e25_blk00000e26_sig000020ba,
      A2 => blk00000e25_blk00000e26_sig000020b9,
      A3 => blk00000e25_blk00000e26_sig000020ba,
      CE => ce,
      CLK => clk,
      D => sig00000cce,
      Q => blk00000e25_blk00000e26_sig000020bf,
      Q15 => NLW_blk00000e25_blk00000e26_blk00000e31_Q15_UNCONNECTED
    );
  blk00000e25_blk00000e26_blk00000e30 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000e25_blk00000e26_sig000020be,
      Q => sig000000c8
    );
  blk00000e25_blk00000e26_blk00000e2f : SRLC16E
    generic map(
      INIT => X"0000"
    )
    port map (
      A0 => blk00000e25_blk00000e26_sig000020b9,
      A1 => blk00000e25_blk00000e26_sig000020ba,
      A2 => blk00000e25_blk00000e26_sig000020b9,
      A3 => blk00000e25_blk00000e26_sig000020ba,
      CE => ce,
      CLK => clk,
      D => sig00000cd0,
      Q => blk00000e25_blk00000e26_sig000020be,
      Q15 => NLW_blk00000e25_blk00000e26_blk00000e2f_Q15_UNCONNECTED
    );
  blk00000e25_blk00000e26_blk00000e2e : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000e25_blk00000e26_sig000020bd,
      Q => sig000000c4
    );
  blk00000e25_blk00000e26_blk00000e2d : SRLC16E
    generic map(
      INIT => X"0000"
    )
    port map (
      A0 => blk00000e25_blk00000e26_sig000020b9,
      A1 => blk00000e25_blk00000e26_sig000020ba,
      A2 => blk00000e25_blk00000e26_sig000020b9,
      A3 => blk00000e25_blk00000e26_sig000020ba,
      CE => ce,
      CLK => clk,
      D => sig00000ccc,
      Q => blk00000e25_blk00000e26_sig000020bd,
      Q15 => NLW_blk00000e25_blk00000e26_blk00000e2d_Q15_UNCONNECTED
    );
  blk00000e25_blk00000e26_blk00000e2c : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000e25_blk00000e26_sig000020bc,
      Q => sig000000c3
    );
  blk00000e25_blk00000e26_blk00000e2b : SRLC16E
    generic map(
      INIT => X"0000"
    )
    port map (
      A0 => blk00000e25_blk00000e26_sig000020b9,
      A1 => blk00000e25_blk00000e26_sig000020ba,
      A2 => blk00000e25_blk00000e26_sig000020b9,
      A3 => blk00000e25_blk00000e26_sig000020ba,
      CE => ce,
      CLK => clk,
      D => sig00000ccb,
      Q => blk00000e25_blk00000e26_sig000020bc,
      Q15 => NLW_blk00000e25_blk00000e26_blk00000e2b_Q15_UNCONNECTED
    );
  blk00000e25_blk00000e26_blk00000e2a : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000e25_blk00000e26_sig000020bb,
      Q => sig000000c5
    );
  blk00000e25_blk00000e26_blk00000e29 : SRLC16E
    generic map(
      INIT => X"0000"
    )
    port map (
      A0 => blk00000e25_blk00000e26_sig000020b9,
      A1 => blk00000e25_blk00000e26_sig000020ba,
      A2 => blk00000e25_blk00000e26_sig000020b9,
      A3 => blk00000e25_blk00000e26_sig000020ba,
      CE => ce,
      CLK => clk,
      D => sig00000ccd,
      Q => blk00000e25_blk00000e26_sig000020bb,
      Q15 => NLW_blk00000e25_blk00000e26_blk00000e29_Q15_UNCONNECTED
    );
  blk00000e25_blk00000e26_blk00000e28 : VCC
    port map (
      P => blk00000e25_blk00000e26_sig000020ba
    );
  blk00000e25_blk00000e26_blk00000e27 : GND
    port map (
      G => blk00000e25_blk00000e26_sig000020b9
    );
  blk00000e35_blk00000e6d : LUT2
    generic map(
      INIT => X"9"
    )
    port map (
      I0 => sig00000e8e,
      I1 => sig00000e64,
      O => blk00000e35_sig000020fe
    );
  blk00000e35_blk00000e6c : LUT2
    generic map(
      INIT => X"9"
    )
    port map (
      I0 => sig00000e8d,
      I1 => sig00000e63,
      O => blk00000e35_sig000020ff
    );
  blk00000e35_blk00000e6b : LUT2
    generic map(
      INIT => X"9"
    )
    port map (
      I0 => sig00000e8c,
      I1 => sig00000e62,
      O => blk00000e35_sig00002100
    );
  blk00000e35_blk00000e6a : LUT2
    generic map(
      INIT => X"9"
    )
    port map (
      I0 => sig00000e8b,
      I1 => sig00000e61,
      O => blk00000e35_sig00002101
    );
  blk00000e35_blk00000e69 : LUT2
    generic map(
      INIT => X"9"
    )
    port map (
      I0 => sig00000e8a,
      I1 => sig00000e60,
      O => blk00000e35_sig00002102
    );
  blk00000e35_blk00000e68 : LUT2
    generic map(
      INIT => X"9"
    )
    port map (
      I0 => sig00000e89,
      I1 => sig00000e5f,
      O => blk00000e35_sig00002103
    );
  blk00000e35_blk00000e67 : LUT2
    generic map(
      INIT => X"9"
    )
    port map (
      I0 => sig00000e88,
      I1 => sig00000e5e,
      O => blk00000e35_sig00002104
    );
  blk00000e35_blk00000e66 : LUT2
    generic map(
      INIT => X"9"
    )
    port map (
      I0 => sig00000e87,
      I1 => sig00000e5d,
      O => blk00000e35_sig00002105
    );
  blk00000e35_blk00000e65 : LUT2
    generic map(
      INIT => X"9"
    )
    port map (
      I0 => sig00000e86,
      I1 => sig00000e5c,
      O => blk00000e35_sig00002106
    );
  blk00000e35_blk00000e64 : LUT2
    generic map(
      INIT => X"9"
    )
    port map (
      I0 => sig00000e92,
      I1 => sig00000e68,
      O => blk00000e35_sig00002107
    );
  blk00000e35_blk00000e63 : LUT2
    generic map(
      INIT => X"9"
    )
    port map (
      I0 => sig00000e91,
      I1 => sig00000e67,
      O => blk00000e35_sig000020fb
    );
  blk00000e35_blk00000e62 : LUT2
    generic map(
      INIT => X"9"
    )
    port map (
      I0 => sig00000e90,
      I1 => sig00000e66,
      O => blk00000e35_sig000020fc
    );
  blk00000e35_blk00000e61 : LUT2
    generic map(
      INIT => X"9"
    )
    port map (
      I0 => sig00000e8f,
      I1 => sig00000e65,
      O => blk00000e35_sig000020fd
    );
  blk00000e35_blk00000e60 : LUT2
    generic map(
      INIT => X"9"
    )
    port map (
      I0 => sig00000e85,
      I1 => sig00000e5b,
      O => blk00000e35_sig00002108
    );
  blk00000e35_blk00000e5f : MUXCY
    port map (
      CI => blk00000e35_sig00002116,
      DI => sig00000e85,
      S => blk00000e35_sig00002108,
      O => blk00000e35_sig00002115
    );
  blk00000e35_blk00000e5e : MUXCY
    port map (
      CI => blk00000e35_sig00002115,
      DI => sig00000e86,
      S => blk00000e35_sig00002106,
      O => blk00000e35_sig00002114
    );
  blk00000e35_blk00000e5d : MUXCY
    port map (
      CI => blk00000e35_sig00002114,
      DI => sig00000e87,
      S => blk00000e35_sig00002105,
      O => blk00000e35_sig00002113
    );
  blk00000e35_blk00000e5c : MUXCY
    port map (
      CI => blk00000e35_sig00002113,
      DI => sig00000e88,
      S => blk00000e35_sig00002104,
      O => blk00000e35_sig00002112
    );
  blk00000e35_blk00000e5b : MUXCY
    port map (
      CI => blk00000e35_sig00002112,
      DI => sig00000e89,
      S => blk00000e35_sig00002103,
      O => blk00000e35_sig00002111
    );
  blk00000e35_blk00000e5a : MUXCY
    port map (
      CI => blk00000e35_sig00002111,
      DI => sig00000e8a,
      S => blk00000e35_sig00002102,
      O => blk00000e35_sig00002110
    );
  blk00000e35_blk00000e59 : MUXCY
    port map (
      CI => blk00000e35_sig00002110,
      DI => sig00000e8b,
      S => blk00000e35_sig00002101,
      O => blk00000e35_sig0000210f
    );
  blk00000e35_blk00000e58 : MUXCY
    port map (
      CI => blk00000e35_sig0000210f,
      DI => sig00000e8c,
      S => blk00000e35_sig00002100,
      O => blk00000e35_sig0000210e
    );
  blk00000e35_blk00000e57 : MUXCY
    port map (
      CI => blk00000e35_sig0000210e,
      DI => sig00000e8d,
      S => blk00000e35_sig000020ff,
      O => blk00000e35_sig0000210d
    );
  blk00000e35_blk00000e56 : MUXCY
    port map (
      CI => blk00000e35_sig0000210d,
      DI => sig00000e8e,
      S => blk00000e35_sig000020fe,
      O => blk00000e35_sig0000210c
    );
  blk00000e35_blk00000e55 : MUXCY
    port map (
      CI => blk00000e35_sig0000210c,
      DI => sig00000e8f,
      S => blk00000e35_sig000020fd,
      O => blk00000e35_sig0000210b
    );
  blk00000e35_blk00000e54 : MUXCY
    port map (
      CI => blk00000e35_sig0000210b,
      DI => sig00000e90,
      S => blk00000e35_sig000020fc,
      O => blk00000e35_sig0000210a
    );
  blk00000e35_blk00000e53 : MUXCY
    port map (
      CI => blk00000e35_sig0000210a,
      DI => sig00000e91,
      S => blk00000e35_sig000020fb,
      O => blk00000e35_sig00002109
    );
  blk00000e35_blk00000e52 : XORCY
    port map (
      CI => blk00000e35_sig00002116,
      LI => blk00000e35_sig00002108,
      O => blk00000e35_sig000020fa
    );
  blk00000e35_blk00000e51 : XORCY
    port map (
      CI => blk00000e35_sig00002115,
      LI => blk00000e35_sig00002106,
      O => blk00000e35_sig000020f9
    );
  blk00000e35_blk00000e50 : XORCY
    port map (
      CI => blk00000e35_sig00002114,
      LI => blk00000e35_sig00002105,
      O => blk00000e35_sig000020f8
    );
  blk00000e35_blk00000e4f : XORCY
    port map (
      CI => blk00000e35_sig00002113,
      LI => blk00000e35_sig00002104,
      O => blk00000e35_sig000020f7
    );
  blk00000e35_blk00000e4e : XORCY
    port map (
      CI => blk00000e35_sig00002112,
      LI => blk00000e35_sig00002103,
      O => blk00000e35_sig000020f6
    );
  blk00000e35_blk00000e4d : XORCY
    port map (
      CI => blk00000e35_sig00002111,
      LI => blk00000e35_sig00002102,
      O => blk00000e35_sig000020f5
    );
  blk00000e35_blk00000e4c : XORCY
    port map (
      CI => blk00000e35_sig00002110,
      LI => blk00000e35_sig00002101,
      O => blk00000e35_sig000020f4
    );
  blk00000e35_blk00000e4b : XORCY
    port map (
      CI => blk00000e35_sig0000210f,
      LI => blk00000e35_sig00002100,
      O => blk00000e35_sig000020f3
    );
  blk00000e35_blk00000e4a : XORCY
    port map (
      CI => blk00000e35_sig0000210e,
      LI => blk00000e35_sig000020ff,
      O => blk00000e35_sig000020f2
    );
  blk00000e35_blk00000e49 : XORCY
    port map (
      CI => blk00000e35_sig0000210d,
      LI => blk00000e35_sig000020fe,
      O => blk00000e35_sig000020f1
    );
  blk00000e35_blk00000e48 : XORCY
    port map (
      CI => blk00000e35_sig0000210c,
      LI => blk00000e35_sig000020fd,
      O => blk00000e35_sig000020f0
    );
  blk00000e35_blk00000e47 : XORCY
    port map (
      CI => blk00000e35_sig0000210b,
      LI => blk00000e35_sig000020fc,
      O => blk00000e35_sig000020ef
    );
  blk00000e35_blk00000e46 : XORCY
    port map (
      CI => blk00000e35_sig0000210a,
      LI => blk00000e35_sig000020fb,
      O => blk00000e35_sig000020ee
    );
  blk00000e35_blk00000e45 : XORCY
    port map (
      CI => blk00000e35_sig00002109,
      LI => blk00000e35_sig00002107,
      O => blk00000e35_sig000020ed
    );
  blk00000e35_blk00000e44 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000e35_sig000020ed,
      Q => sig00000e4c
    );
  blk00000e35_blk00000e43 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000e35_sig000020ee,
      Q => sig00000e4b
    );
  blk00000e35_blk00000e42 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000e35_sig000020ef,
      Q => sig00000e4a
    );
  blk00000e35_blk00000e41 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000e35_sig000020f0,
      Q => sig00000e49
    );
  blk00000e35_blk00000e40 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000e35_sig000020f1,
      Q => sig00000e48
    );
  blk00000e35_blk00000e3f : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000e35_sig000020f2,
      Q => sig00000e47
    );
  blk00000e35_blk00000e3e : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000e35_sig000020f3,
      Q => sig00000e46
    );
  blk00000e35_blk00000e3d : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000e35_sig000020f4,
      Q => sig00000e45
    );
  blk00000e35_blk00000e3c : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000e35_sig000020f5,
      Q => sig00000e44
    );
  blk00000e35_blk00000e3b : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000e35_sig000020f6,
      Q => sig00000e43
    );
  blk00000e35_blk00000e3a : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000e35_sig000020f7,
      Q => sig00000e42
    );
  blk00000e35_blk00000e39 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000e35_sig000020f8,
      Q => sig00000e41
    );
  blk00000e35_blk00000e38 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000e35_sig000020f9,
      Q => sig00000e40
    );
  blk00000e35_blk00000e37 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000e35_sig000020fa,
      Q => sig00000e3f
    );
  blk00000e35_blk00000e36 : VCC
    port map (
      P => blk00000e35_sig00002116
    );
  blk00000e6e_blk00000ea6 : LUT2
    generic map(
      INIT => X"6"
    )
    port map (
      I0 => sig00000e8e,
      I1 => sig00000e64,
      O => blk00000e6e_sig00002155
    );
  blk00000e6e_blk00000ea5 : LUT2
    generic map(
      INIT => X"6"
    )
    port map (
      I0 => sig00000e8d,
      I1 => sig00000e63,
      O => blk00000e6e_sig00002156
    );
  blk00000e6e_blk00000ea4 : LUT2
    generic map(
      INIT => X"6"
    )
    port map (
      I0 => sig00000e8c,
      I1 => sig00000e62,
      O => blk00000e6e_sig00002157
    );
  blk00000e6e_blk00000ea3 : LUT2
    generic map(
      INIT => X"6"
    )
    port map (
      I0 => sig00000e8b,
      I1 => sig00000e61,
      O => blk00000e6e_sig00002158
    );
  blk00000e6e_blk00000ea2 : LUT2
    generic map(
      INIT => X"6"
    )
    port map (
      I0 => sig00000e8a,
      I1 => sig00000e60,
      O => blk00000e6e_sig00002159
    );
  blk00000e6e_blk00000ea1 : LUT2
    generic map(
      INIT => X"6"
    )
    port map (
      I0 => sig00000e89,
      I1 => sig00000e5f,
      O => blk00000e6e_sig0000215a
    );
  blk00000e6e_blk00000ea0 : LUT2
    generic map(
      INIT => X"6"
    )
    port map (
      I0 => sig00000e88,
      I1 => sig00000e5e,
      O => blk00000e6e_sig0000215b
    );
  blk00000e6e_blk00000e9f : LUT2
    generic map(
      INIT => X"6"
    )
    port map (
      I0 => sig00000e87,
      I1 => sig00000e5d,
      O => blk00000e6e_sig0000215c
    );
  blk00000e6e_blk00000e9e : LUT2
    generic map(
      INIT => X"6"
    )
    port map (
      I0 => sig00000e86,
      I1 => sig00000e5c,
      O => blk00000e6e_sig0000215d
    );
  blk00000e6e_blk00000e9d : LUT2
    generic map(
      INIT => X"6"
    )
    port map (
      I0 => sig00000e92,
      I1 => sig00000e68,
      O => blk00000e6e_sig0000215e
    );
  blk00000e6e_blk00000e9c : LUT2
    generic map(
      INIT => X"6"
    )
    port map (
      I0 => sig00000e91,
      I1 => sig00000e67,
      O => blk00000e6e_sig00002152
    );
  blk00000e6e_blk00000e9b : LUT2
    generic map(
      INIT => X"6"
    )
    port map (
      I0 => sig00000e90,
      I1 => sig00000e66,
      O => blk00000e6e_sig00002153
    );
  blk00000e6e_blk00000e9a : LUT2
    generic map(
      INIT => X"6"
    )
    port map (
      I0 => sig00000e8f,
      I1 => sig00000e65,
      O => blk00000e6e_sig00002154
    );
  blk00000e6e_blk00000e99 : LUT2
    generic map(
      INIT => X"6"
    )
    port map (
      I0 => sig00000e85,
      I1 => sig00000e5b,
      O => blk00000e6e_sig0000215f
    );
  blk00000e6e_blk00000e98 : MUXCY
    port map (
      CI => blk00000e6e_sig00002143,
      DI => sig00000e85,
      S => blk00000e6e_sig0000215f,
      O => blk00000e6e_sig0000216c
    );
  blk00000e6e_blk00000e97 : MUXCY
    port map (
      CI => blk00000e6e_sig0000216c,
      DI => sig00000e86,
      S => blk00000e6e_sig0000215d,
      O => blk00000e6e_sig0000216b
    );
  blk00000e6e_blk00000e96 : MUXCY
    port map (
      CI => blk00000e6e_sig0000216b,
      DI => sig00000e87,
      S => blk00000e6e_sig0000215c,
      O => blk00000e6e_sig0000216a
    );
  blk00000e6e_blk00000e95 : MUXCY
    port map (
      CI => blk00000e6e_sig0000216a,
      DI => sig00000e88,
      S => blk00000e6e_sig0000215b,
      O => blk00000e6e_sig00002169
    );
  blk00000e6e_blk00000e94 : MUXCY
    port map (
      CI => blk00000e6e_sig00002169,
      DI => sig00000e89,
      S => blk00000e6e_sig0000215a,
      O => blk00000e6e_sig00002168
    );
  blk00000e6e_blk00000e93 : MUXCY
    port map (
      CI => blk00000e6e_sig00002168,
      DI => sig00000e8a,
      S => blk00000e6e_sig00002159,
      O => blk00000e6e_sig00002167
    );
  blk00000e6e_blk00000e92 : MUXCY
    port map (
      CI => blk00000e6e_sig00002167,
      DI => sig00000e8b,
      S => blk00000e6e_sig00002158,
      O => blk00000e6e_sig00002166
    );
  blk00000e6e_blk00000e91 : MUXCY
    port map (
      CI => blk00000e6e_sig00002166,
      DI => sig00000e8c,
      S => blk00000e6e_sig00002157,
      O => blk00000e6e_sig00002165
    );
  blk00000e6e_blk00000e90 : MUXCY
    port map (
      CI => blk00000e6e_sig00002165,
      DI => sig00000e8d,
      S => blk00000e6e_sig00002156,
      O => blk00000e6e_sig00002164
    );
  blk00000e6e_blk00000e8f : MUXCY
    port map (
      CI => blk00000e6e_sig00002164,
      DI => sig00000e8e,
      S => blk00000e6e_sig00002155,
      O => blk00000e6e_sig00002163
    );
  blk00000e6e_blk00000e8e : MUXCY
    port map (
      CI => blk00000e6e_sig00002163,
      DI => sig00000e8f,
      S => blk00000e6e_sig00002154,
      O => blk00000e6e_sig00002162
    );
  blk00000e6e_blk00000e8d : MUXCY
    port map (
      CI => blk00000e6e_sig00002162,
      DI => sig00000e90,
      S => blk00000e6e_sig00002153,
      O => blk00000e6e_sig00002161
    );
  blk00000e6e_blk00000e8c : MUXCY
    port map (
      CI => blk00000e6e_sig00002161,
      DI => sig00000e91,
      S => blk00000e6e_sig00002152,
      O => blk00000e6e_sig00002160
    );
  blk00000e6e_blk00000e8b : XORCY
    port map (
      CI => blk00000e6e_sig00002143,
      LI => blk00000e6e_sig0000215f,
      O => blk00000e6e_sig00002151
    );
  blk00000e6e_blk00000e8a : XORCY
    port map (
      CI => blk00000e6e_sig0000216c,
      LI => blk00000e6e_sig0000215d,
      O => blk00000e6e_sig00002150
    );
  blk00000e6e_blk00000e89 : XORCY
    port map (
      CI => blk00000e6e_sig0000216b,
      LI => blk00000e6e_sig0000215c,
      O => blk00000e6e_sig0000214f
    );
  blk00000e6e_blk00000e88 : XORCY
    port map (
      CI => blk00000e6e_sig0000216a,
      LI => blk00000e6e_sig0000215b,
      O => blk00000e6e_sig0000214e
    );
  blk00000e6e_blk00000e87 : XORCY
    port map (
      CI => blk00000e6e_sig00002169,
      LI => blk00000e6e_sig0000215a,
      O => blk00000e6e_sig0000214d
    );
  blk00000e6e_blk00000e86 : XORCY
    port map (
      CI => blk00000e6e_sig00002168,
      LI => blk00000e6e_sig00002159,
      O => blk00000e6e_sig0000214c
    );
  blk00000e6e_blk00000e85 : XORCY
    port map (
      CI => blk00000e6e_sig00002167,
      LI => blk00000e6e_sig00002158,
      O => blk00000e6e_sig0000214b
    );
  blk00000e6e_blk00000e84 : XORCY
    port map (
      CI => blk00000e6e_sig00002166,
      LI => blk00000e6e_sig00002157,
      O => blk00000e6e_sig0000214a
    );
  blk00000e6e_blk00000e83 : XORCY
    port map (
      CI => blk00000e6e_sig00002165,
      LI => blk00000e6e_sig00002156,
      O => blk00000e6e_sig00002149
    );
  blk00000e6e_blk00000e82 : XORCY
    port map (
      CI => blk00000e6e_sig00002164,
      LI => blk00000e6e_sig00002155,
      O => blk00000e6e_sig00002148
    );
  blk00000e6e_blk00000e81 : XORCY
    port map (
      CI => blk00000e6e_sig00002163,
      LI => blk00000e6e_sig00002154,
      O => blk00000e6e_sig00002147
    );
  blk00000e6e_blk00000e80 : XORCY
    port map (
      CI => blk00000e6e_sig00002162,
      LI => blk00000e6e_sig00002153,
      O => blk00000e6e_sig00002146
    );
  blk00000e6e_blk00000e7f : XORCY
    port map (
      CI => blk00000e6e_sig00002161,
      LI => blk00000e6e_sig00002152,
      O => blk00000e6e_sig00002145
    );
  blk00000e6e_blk00000e7e : XORCY
    port map (
      CI => blk00000e6e_sig00002160,
      LI => blk00000e6e_sig0000215e,
      O => blk00000e6e_sig00002144
    );
  blk00000e6e_blk00000e7d : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000e6e_sig00002144,
      Q => sig00000e5a
    );
  blk00000e6e_blk00000e7c : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000e6e_sig00002145,
      Q => sig00000e59
    );
  blk00000e6e_blk00000e7b : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000e6e_sig00002146,
      Q => sig00000e58
    );
  blk00000e6e_blk00000e7a : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000e6e_sig00002147,
      Q => sig00000e57
    );
  blk00000e6e_blk00000e79 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000e6e_sig00002148,
      Q => sig00000e56
    );
  blk00000e6e_blk00000e78 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000e6e_sig00002149,
      Q => sig00000e55
    );
  blk00000e6e_blk00000e77 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000e6e_sig0000214a,
      Q => sig00000e54
    );
  blk00000e6e_blk00000e76 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000e6e_sig0000214b,
      Q => sig00000e53
    );
  blk00000e6e_blk00000e75 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000e6e_sig0000214c,
      Q => sig00000e52
    );
  blk00000e6e_blk00000e74 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000e6e_sig0000214d,
      Q => sig00000e51
    );
  blk00000e6e_blk00000e73 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000e6e_sig0000214e,
      Q => sig00000e50
    );
  blk00000e6e_blk00000e72 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000e6e_sig0000214f,
      Q => sig00000e4f
    );
  blk00000e6e_blk00000e71 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000e6e_sig00002150,
      Q => sig00000e4e
    );
  blk00000e6e_blk00000e70 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000e6e_sig00002151,
      Q => sig00000e4d
    );
  blk00000e6e_blk00000e6f : GND
    port map (
      G => blk00000e6e_sig00002143
    );
  blk00000ea7_blk00000ea8_blk00000eab : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000ea7_blk00000ea8_sig0000217d,
      Q => sig00000eb1
    );
  blk00000ea7_blk00000ea8_blk00000eaa : SRLC16E
    generic map(
      INIT => X"0000"
    )
    port map (
      A0 => blk00000ea7_blk00000ea8_sig0000217c,
      A1 => blk00000ea7_blk00000ea8_sig0000217c,
      A2 => blk00000ea7_blk00000ea8_sig0000217c,
      A3 => blk00000ea7_blk00000ea8_sig0000217c,
      CE => ce,
      CLK => clk,
      D => sig00000eb2,
      Q => blk00000ea7_blk00000ea8_sig0000217d,
      Q15 => NLW_blk00000ea7_blk00000ea8_blk00000eaa_Q15_UNCONNECTED
    );
  blk00000ea7_blk00000ea8_blk00000ea9 : GND
    port map (
      G => blk00000ea7_blk00000ea8_sig0000217c
    );
  blk00000eac_blk00000ead_blk00000eb0 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000eac_blk00000ead_sig0000218e,
      Q => sig00000eb2
    );
  blk00000eac_blk00000ead_blk00000eaf : SRLC16E
    generic map(
      INIT => X"0000"
    )
    port map (
      A0 => blk00000eac_blk00000ead_sig0000218d,
      A1 => blk00000eac_blk00000ead_sig0000218d,
      A2 => blk00000eac_blk00000ead_sig0000218d,
      A3 => blk00000eac_blk00000ead_sig0000218d,
      CE => ce,
      CLK => clk,
      D => sig00000eb3,
      Q => blk00000eac_blk00000ead_sig0000218e,
      Q15 => NLW_blk00000eac_blk00000ead_blk00000eaf_Q15_UNCONNECTED
    );
  blk00000eac_blk00000ead_blk00000eae : GND
    port map (
      G => blk00000eac_blk00000ead_sig0000218d
    );
  blk00000fbf_blk00000fc1 : RAMB18SDP
    generic map(
      DO_REG => 1,
      INIT => X"000000000",
      INITP_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INITP_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INITP_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INITP_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INITP_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INITP_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INITP_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INITP_07 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_07 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_08 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_09 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_0F => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_10 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_11 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_12 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_13 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_14 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_15 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_16 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_17 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_18 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_19 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_1A => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_1B => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_1C => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_1D => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_1E => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_1F => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_20 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_21 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_22 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_23 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_24 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_25 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_26 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_27 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_28 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_29 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_2A => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_2B => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_2C => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_2D => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_2E => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_2F => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_30 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_31 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_32 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_33 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_34 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_FILE => "NONE",
      SIM_COLLISION_CHECK => "GENERATE_X_ONLY",
      SIM_MODE => "SAFE",
      SRVAL => X"000000000"
    )
    port map (
      RDCLK => clk,
      WRCLK => clk,
      RDEN => ce,
      WREN => ce,
      REGCE => ce,
      SSR => blk00000fbf_sig000021cf,
      RDADDR(8) => sig00000057,
      RDADDR(7) => sig00000056,
      RDADDR(6) => sig00000055,
      RDADDR(5) => sig00000054,
      RDADDR(4) => sig00000053,
      RDADDR(3) => sig00000052,
      RDADDR(2) => blk00000fbf_sig000021cf,
      RDADDR(1) => blk00000fbf_sig000021cf,
      RDADDR(0) => blk00000fbf_sig000021cf,
      WRADDR(8) => sig0000005d,
      WRADDR(7) => sig0000005c,
      WRADDR(6) => sig0000005b,
      WRADDR(5) => sig0000005a,
      WRADDR(4) => sig00000059,
      WRADDR(3) => sig00000058,
      WRADDR(2) => blk00000fbf_sig000021cf,
      WRADDR(1) => blk00000fbf_sig000021cf,
      WRADDR(0) => blk00000fbf_sig000021cf,
      DI(31) => blk00000fbf_sig000021cf,
      DI(30) => blk00000fbf_sig000021cf,
      DI(29) => blk00000fbf_sig000021cf,
      DI(28) => blk00000fbf_sig000021cf,
      DI(27) => blk00000fbf_sig000021cf,
      DI(26) => blk00000fbf_sig000021cf,
      DI(25) => blk00000fbf_sig000021cf,
      DI(24) => blk00000fbf_sig000021cf,
      DI(23) => blk00000fbf_sig000021cf,
      DI(22) => blk00000fbf_sig000021cf,
      DI(21) => sig00000092,
      DI(20) => sig00000091,
      DI(19) => sig00000090,
      DI(18) => sig0000008f,
      DI(17) => sig0000008e,
      DI(16) => sig0000008d,
      DI(15) => sig0000008b,
      DI(14) => sig0000008a,
      DI(13) => sig00000089,
      DI(12) => sig00000088,
      DI(11) => sig00000087,
      DI(10) => sig00000086,
      DI(9) => sig00000085,
      DI(8) => sig00000084,
      DI(7) => sig00000082,
      DI(6) => sig00000081,
      DI(5) => sig00000080,
      DI(4) => sig0000007f,
      DI(3) => sig0000007e,
      DI(2) => sig0000007d,
      DI(1) => sig0000007c,
      DI(0) => sig0000007b,
      DIP(3) => blk00000fbf_sig000021cf,
      DIP(2) => blk00000fbf_sig000021cf,
      DIP(1) => sig0000008c,
      DIP(0) => sig00000083,
      DO(31) => NLW_blk00000fbf_blk00000fc1_DO_31_UNCONNECTED,
      DO(30) => NLW_blk00000fbf_blk00000fc1_DO_30_UNCONNECTED,
      DO(29) => NLW_blk00000fbf_blk00000fc1_DO_29_UNCONNECTED,
      DO(28) => NLW_blk00000fbf_blk00000fc1_DO_28_UNCONNECTED,
      DO(27) => NLW_blk00000fbf_blk00000fc1_DO_27_UNCONNECTED,
      DO(26) => NLW_blk00000fbf_blk00000fc1_DO_26_UNCONNECTED,
      DO(25) => NLW_blk00000fbf_blk00000fc1_DO_25_UNCONNECTED,
      DO(24) => NLW_blk00000fbf_blk00000fc1_DO_24_UNCONNECTED,
      DO(23) => NLW_blk00000fbf_blk00000fc1_DO_23_UNCONNECTED,
      DO(22) => NLW_blk00000fbf_blk00000fc1_DO_22_UNCONNECTED,
      DO(21) => sig0000007a,
      DO(20) => sig00000079,
      DO(19) => sig00000078,
      DO(18) => sig00000077,
      DO(17) => sig00000076,
      DO(16) => sig00000075,
      DO(15) => sig00000073,
      DO(14) => sig00000072,
      DO(13) => sig00000071,
      DO(12) => sig00000070,
      DO(11) => sig0000006f,
      DO(10) => sig0000006e,
      DO(9) => sig0000006d,
      DO(8) => sig0000006c,
      DO(7) => sig0000006a,
      DO(6) => sig00000069,
      DO(5) => sig00000068,
      DO(4) => sig00000067,
      DO(3) => sig00000066,
      DO(2) => sig00000065,
      DO(1) => sig00000064,
      DO(0) => sig00000063,
      DOP(3) => NLW_blk00000fbf_blk00000fc1_DOP_3_UNCONNECTED,
      DOP(2) => NLW_blk00000fbf_blk00000fc1_DOP_2_UNCONNECTED,
      DOP(1) => sig00000074,
      DOP(0) => sig0000006b,
      WE(3) => sig000000a1,
      WE(2) => sig000000a1,
      WE(1) => sig000000a1,
      WE(0) => sig000000a1
    );
  blk00000fbf_blk00000fc0 : GND
    port map (
      G => blk00000fbf_sig000021cf
    );
  blk00000fc2_blk00000fc3_blk00000fd1 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000fc2_blk00000fc3_sig000021f4,
      Q => sig00000ee1
    );
  blk00000fc2_blk00000fc3_blk00000fd0 : SRLC16E
    generic map(
      INIT => X"0000"
    )
    port map (
      A0 => blk00000fc2_blk00000fc3_sig000021ee,
      A1 => blk00000fc2_blk00000fc3_sig000021ed,
      A2 => blk00000fc2_blk00000fc3_sig000021ed,
      A3 => blk00000fc2_blk00000fc3_sig000021ed,
      CE => ce,
      CLK => clk,
      D => sig0000009f,
      Q => blk00000fc2_blk00000fc3_sig000021f4,
      Q15 => NLW_blk00000fc2_blk00000fc3_blk00000fd0_Q15_UNCONNECTED
    );
  blk00000fc2_blk00000fc3_blk00000fcf : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000fc2_blk00000fc3_sig000021f3,
      Q => sig00000ee0
    );
  blk00000fc2_blk00000fc3_blk00000fce : SRLC16E
    generic map(
      INIT => X"0000"
    )
    port map (
      A0 => blk00000fc2_blk00000fc3_sig000021ee,
      A1 => blk00000fc2_blk00000fc3_sig000021ed,
      A2 => blk00000fc2_blk00000fc3_sig000021ed,
      A3 => blk00000fc2_blk00000fc3_sig000021ed,
      CE => ce,
      CLK => clk,
      D => sig0000009e,
      Q => blk00000fc2_blk00000fc3_sig000021f3,
      Q15 => NLW_blk00000fc2_blk00000fc3_blk00000fce_Q15_UNCONNECTED
    );
  blk00000fc2_blk00000fc3_blk00000fcd : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000fc2_blk00000fc3_sig000021f2,
      Q => sig00000ee2
    );
  blk00000fc2_blk00000fc3_blk00000fcc : SRLC16E
    generic map(
      INIT => X"0000"
    )
    port map (
      A0 => blk00000fc2_blk00000fc3_sig000021ee,
      A1 => blk00000fc2_blk00000fc3_sig000021ed,
      A2 => blk00000fc2_blk00000fc3_sig000021ed,
      A3 => blk00000fc2_blk00000fc3_sig000021ed,
      CE => ce,
      CLK => clk,
      D => sig000000a0,
      Q => blk00000fc2_blk00000fc3_sig000021f2,
      Q15 => NLW_blk00000fc2_blk00000fc3_blk00000fcc_Q15_UNCONNECTED
    );
  blk00000fc2_blk00000fc3_blk00000fcb : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000fc2_blk00000fc3_sig000021f1,
      Q => sig00000ede
    );
  blk00000fc2_blk00000fc3_blk00000fca : SRLC16E
    generic map(
      INIT => X"0000"
    )
    port map (
      A0 => blk00000fc2_blk00000fc3_sig000021ee,
      A1 => blk00000fc2_blk00000fc3_sig000021ed,
      A2 => blk00000fc2_blk00000fc3_sig000021ed,
      A3 => blk00000fc2_blk00000fc3_sig000021ed,
      CE => ce,
      CLK => clk,
      D => sig0000009c,
      Q => blk00000fc2_blk00000fc3_sig000021f1,
      Q15 => NLW_blk00000fc2_blk00000fc3_blk00000fca_Q15_UNCONNECTED
    );
  blk00000fc2_blk00000fc3_blk00000fc9 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000fc2_blk00000fc3_sig000021f0,
      Q => sig00000edd
    );
  blk00000fc2_blk00000fc3_blk00000fc8 : SRLC16E
    generic map(
      INIT => X"0000"
    )
    port map (
      A0 => blk00000fc2_blk00000fc3_sig000021ee,
      A1 => blk00000fc2_blk00000fc3_sig000021ed,
      A2 => blk00000fc2_blk00000fc3_sig000021ed,
      A3 => blk00000fc2_blk00000fc3_sig000021ed,
      CE => ce,
      CLK => clk,
      D => sig0000009b,
      Q => blk00000fc2_blk00000fc3_sig000021f0,
      Q15 => NLW_blk00000fc2_blk00000fc3_blk00000fc8_Q15_UNCONNECTED
    );
  blk00000fc2_blk00000fc3_blk00000fc7 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000fc2_blk00000fc3_sig000021ef,
      Q => sig00000edf
    );
  blk00000fc2_blk00000fc3_blk00000fc6 : SRLC16E
    generic map(
      INIT => X"0000"
    )
    port map (
      A0 => blk00000fc2_blk00000fc3_sig000021ee,
      A1 => blk00000fc2_blk00000fc3_sig000021ed,
      A2 => blk00000fc2_blk00000fc3_sig000021ed,
      A3 => blk00000fc2_blk00000fc3_sig000021ed,
      CE => ce,
      CLK => clk,
      D => sig0000009d,
      Q => blk00000fc2_blk00000fc3_sig000021ef,
      Q15 => NLW_blk00000fc2_blk00000fc3_blk00000fc6_Q15_UNCONNECTED
    );
  blk00000fc2_blk00000fc3_blk00000fc5 : VCC
    port map (
      P => blk00000fc2_blk00000fc3_sig000021ee
    );
  blk00000fc2_blk00000fc3_blk00000fc4 : GND
    port map (
      G => blk00000fc2_blk00000fc3_sig000021ed
    );
  blk00000fd8_blk00000fd9_blk00000fdc : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000fd8_blk00000fd9_sig00002205,
      Q => sig00000ee6
    );
  blk00000fd8_blk00000fd9_blk00000fdb : SRLC16E
    generic map(
      INIT => X"0000"
    )
    port map (
      A0 => blk00000fd8_blk00000fd9_sig00002204,
      A1 => blk00000fd8_blk00000fd9_sig00002204,
      A2 => blk00000fd8_blk00000fd9_sig00002204,
      A3 => blk00000fd8_blk00000fd9_sig00002204,
      CE => ce,
      CLK => clk,
      D => sig0000011d,
      Q => blk00000fd8_blk00000fd9_sig00002205,
      Q15 => NLW_blk00000fd8_blk00000fd9_blk00000fdb_Q15_UNCONNECTED
    );
  blk00000fd8_blk00000fd9_blk00000fda : GND
    port map (
      G => blk00000fd8_blk00000fd9_sig00002204
    );

end STRUCTURE;
