/*
======================================================================================
				Standard   : WIFI
				Block name : BPSK deMapper
======================================================================================
*/
//====================================================================================
module demapper_bpskMod_wifi
(
	clk,
	reset,
	valid_in,
	data_in_real,
	data_in_imag,
	data_out,
	valid_out
);
	//============================================================================	
	input clk;
	input reset;
	input valid_in;
	input [11:0] data_in_real;
	input [11:0] data_in_imag;
	output data_out;
	output valid_out;
	//============================================================================	
	reg valid_out_1;
	reg data_out;
	//============================================================================	
	always@(posedge clk or negedge reset)
	begin
		//====================================================================
		if(!reset)
		begin
			data_out	 	<= 0;
			valid_out_1 	<= 0;
		end
		//====================================================================
		else
		begin
			//============================================================
			if (valid_in)
			begin
				if ($signed(data_in_real[11 -: 9]) < 0)
				begin
					data_out		<= 0;
					valid_out_1 	<= 1;
				end			 
				else if ($signed(data_in_real[11 -: 9]) >= 0)
				begin
					data_out		<= 1;
					valid_out_1 	<= 1;
				end			 
			end
			//============================================================
			else
			begin
				data_out		<= 0;
				valid_out_1 	<= 0;
			end
			//============================================================
		end
		//====================================================================
	end
	//============================================================================
	assign valid_out = valid_out_1;
	//============================================================================
endmodule