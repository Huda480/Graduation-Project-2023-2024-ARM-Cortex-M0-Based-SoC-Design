/////////////////////////////////////////////////////////////////////
////  AHB DMA not mux                                            ////
////                                                             ////
////  Author: Ibrahim Hossam                                     ////
/////////////////////////////////////////////////////////////////////
module not_mux #(
//==========================================================================
// Parameters
//==========================================================================
parameter width = 5)(
//==========================================================================
// Inputs & Outputs
//==========================================================================
input        [width-1:0]    data_in,
input        [width-1:0]    data_in_2,
input                       selector,
output reg   [width-1:0]    data_out
);
//==========================================================================
// Main code
//==========================================================================
    always_comb
    begin
        if(selector)
        data_out = data_in;
        else
        data_out = data_in_2;
    end

endmodule