/////////////////////////////////////////////////////////////////////
////  AHB DMA address increment                                  ////
////                                                             ////
////  Author: Ibrahim Hossam                                     ////
/////////////////////////////////////////////////////////////////////
module ahb_dma_inc30r(
clk,
in,
size_of_incr,
out);
//==========================================================================
// Parameters
//==========================================================================
localparam	INC30_CENTER = 16;
//==========================================================================
// Inputs & Outputs
//==========================================================================
input		clk;
input	[31:0]	in;
input   [2:0]   size_of_incr;
output	[31:0]	out;
//==========================================================================
// Internal signls
//==========================================================================
	reg	[INC30_CENTER:0]	out_r;
//==========================================================================
// Main code
//==========================================================================
	always_comb
	begin
		out_r = in[(INC30_CENTER - 1):0] + (3'b1 << size_of_incr);
	end

	assign out[31:INC30_CENTER] = in[31:INC30_CENTER] + out_r[INC30_CENTER];
	assign out[(INC30_CENTER - 1):0]  = out_r;
endmodule