/*
=====================================================================================
                            Standard    :   All
                            Block name  :   General Clk Distrubution Network  
=====================================================================================
*/
//===================================================================================
`define wifi
//===================================================================================
module clk_distribute
(
    reset,
	clk_200_MHz,
	clk_55_MHz,
	clk_15_MHz,
	clk_100_MHz,
    clk_50_MHz,
    clk_20_MHz_WIFI,
    clk_20_MHz_4G,
    clk_6945_KHz,
    clk_3840_KHz,
    clk_3472_KHz,
    clk_960_KHz,
    clk_480_KHz,
    clk_312_KHz,
    clk_156_KHz
);
	//===============================================================================
	input wire reset;
	input wire clk_200_MHz;
	input wire clk_55_MHz;
	input wire clk_15_MHz;
	output reg clk_100_MHz;
	output reg clk_50_MHz;
	output reg clk_20_MHz_WIFI;
	output reg clk_20_MHz_4G;
	output reg clk_6945_KHz;
	output reg clk_3840_KHz;
	output reg clk_3472_KHz;
	output reg clk_960_KHz;
	output reg clk_480_KHz;
	output reg clk_312_KHz;
    output reg clk_156_KHz;
	//===============================================================================
	reg [1:0] counter_50_MHz;
	reg [2:0] counter_20_MHz_WIFI;
	reg [3:0] counter_20_MHz_4G;
	reg [15:0] counter_312_KHz;
	reg [15:0] counter_156_KHz;
	reg [3:0] divide_8;
	reg [7:0] divide_16;
	reg [15:0] div_32;
    reg [7:0] div_16;
    reg [1:0] div_4;
	//===================================================================================
    `ifdef bluetooth
    //===================================================================================
        always @(posedge clk_55_MHz or negedge reset)
        begin
            //===========================================================================
            if(!reset)
            begin
                clk_6945_KHz            <= 0;
                clk_3472_KHz            <= 0;
                divide_8                <= 0;
                divide_16               <= 0;
            end
            //===========================================================================
            else
            begin
                divide_8[3:0]           <= {divide_8[2:0],!divide_8[3]};        // Dividing by 8
                divide_16[7:0]          <= {divide_16[6:0],!divide_16[7]};      // Dividing by 16 
                clk_6945_KHz            <= !divide_8[3];       
                clk_3472_KHz            <= !divide_16[7];    
            end
            //===========================================================================
        end
    //===================================================================================   
    `elsif three_g
    //===================================================================================
        always @(posedge clk_15_MHz or negedge reset) 
        begin
            //===========================================================================
            if(!reset)
            begin
                clk_3840_KHz            <= 0;
                clk_960_KHz             <= 0;
                clk_480_KHz             <= 0;
                div_32                  <= 0;
                div_16                  <= 0;
                div_4                   <= 0;                  
            end
            //===========================================================================        
            else
            begin
                div_4[1:0]              <= {div_4[0],!div_4[1]} ;            // Dividing by 4
                div_16[7:0]             <= {div_16[6:0],!div_16[7]};        // Dividing by 16
                div_32[15:0]            <= {div_32[14:0],!div_32[15]};      // Dividing by 32
                clk_3840_KHz            <= !div_4[1]; 
                clk_960_KHz             <= !div_16[7];       
                clk_480_KHz             <= !div_32[15];
            end
            //===========================================================================
        end
    //===================================================================================
    `else
    //===================================================================================    	
	always @(posedge clk_200_MHz or negedge reset)
	begin
        //===========================================================================
		if(!reset)
		begin
			clk_100_MHz	             <= 0;
			clk_50_MHz               <= 0;
			clk_20_MHz_WIFI          <= 0;
			clk_20_MHz_4G            <= 0;
			clk_312_KHz	             <= 0;
			clk_156_KHz              <= 0;  
			counter_50_MHz           <= 0;
			counter_20_MHz_WIFI      <= 0;
			counter_20_MHz_4G        <= 0;
			counter_312_KHz          <= 0;
			counter_156_KHz          <= 0;
		end
		//===========================================================================
		else
		begin
            //========================================================================
            `ifdef wifi
            //========================================================================
                clk_100_MHz              <= ~clk_100_MHz;                          // 10 ns
            
                if((counter_50_MHz == 0) | (counter_50_MHz == 2))		          // 20 ns	
				    clk_50_MHz           <= ~clk_50_MHz;
				    
			    if((counter_20_MHz_WIFI == 0) | (counter_20_MHz_WIFI == 5))		  // 25 - 15 ns
				    clk_20_MHz_WIFI      <= ~clk_20_MHz_WIFI;
                
                counter_50_MHz           <= counter_50_MHz + 1;
                counter_20_MHz_WIFI      <= counter_20_MHz_WIFI + 1;
            //========================================================================
            `elsif four_g
            //========================================================================
                if((counter_50_MHz == 0) | (counter_50_MHz == 2))		          // 20 ns	
                    clk_50_MHz           <= ~clk_50_MHz;
                
                if((counter_20_MHz_4G == 0) | (counter_20_MHz_4G == 5))          // 25 - 25 ns
                    clk_20_MHz_4G        <=~ clk_20_MHz_4G;
                    
                counter_20_MHz_4G        <= counter_20_MHz_4G + 1; 
                counter_50_MHz           <= counter_50_MHz + 1;
			    
			    if(counter_20_MHz_4G == 9)
			        counter_20_MHz_4G    <= 0;
            //========================================================================
            `elsif two_g
            //========================================================================
                if((counter_312_KHz == 0) | (counter_312_KHz == 320))            // 3200 ns
                    clk_312_KHz          <= ~clk_312_KHz;
                        
                if((counter_156_KHz == 0) | (counter_156_KHz == 640))           // 6400 ns
                    clk_156_KHz      <= ~clk_156_KHz;            

                counter_312_KHz          <= counter_312_KHz + 1; 
                counter_156_KHz          <= counter_156_KHz + 1;

                if(counter_312_KHz == 639)
                    counter_312_KHz      <= 0;
                
                if(counter_156_KHz == 1279)
                    counter_156_KHz      <= 0;
            //========================================================================
            `else
            `endif
            //========================================================================
		end
		//===========================================================================
	end
	//===============================================================================
	`endif
    //===============================================================================
endmodule