//==============================================================================
// Purpose: SPI Master pkg
// Used in: spi_master
//==============================================================================
package spi_pkg;
  //============================================================================
    //Include new data types
  //============================================================================
      typedef enum logic [1:0] {
          IDLE         = 2'b00,
          CONFIGURE    = 2'b01,
          TRANSFER     = 2'b11,
          TRANSFER_END = 2'b10
      } state_t;
  //============================================================================
endpackage: spi_pkg