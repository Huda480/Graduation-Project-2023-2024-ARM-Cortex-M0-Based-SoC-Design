/////////////////////////////////////////////////////////////////////
////  AHB DMA Definitions                                        ////
////                                                             ////
////  Author: Ibrahim Hossam                                     ////
/////////////////////////////////////////////////////////////////////

`timescale 1ns / 10ps


// CSR Bits
`define	WDMA_CH_EN		0
`define	WDMA_DST_SEL	1
`define	WDMA_SRC_SEL	2
`define	WDMA_INC_DST	3
`define	WDMA_INC_SRC	4
`define	WDMA_MODE		5
`define	WDMA_ARS		6
`define WDMA_USE_ED		7
`define WDMA_WRB		8
`define	WDMA_STOP		9
`define	WDMA_BUSY		10
`define	WDMA_DONE		11
`define	WDMA_ERR		12
`define WDMA_ED_EOL		20

