//===========================================================
// Purpose: Generic Mux select between DIM signals to get only
//          one signal
// Used in: Transpose_mem
//===========================================================
module muxN
#(
    parameter WIDTH = 16,            
    parameter DIM = 8,               
    parameter SEL_WIDTH = $clog2(DIM) 
)
(
    //=======================================================
    // Controls
    //=======================================================
    input  logic        [SEL_WIDTH-1:0] sel_in       ,  
    //=======================================================
    // Inputs    
    //=======================================================
    input  wire logic signed [    WIDTH-1:0] in      [DIM],  
    //=======================================================
    // Outputs
    //=======================================================
    output      logic signed [    WIDTH-1:0] mux_out     
);
    //=======================================================
    // Selection Processs
    //=======================================================
    assign mux_out = in[sel_in];
    //=======================================================
endmodule
