//==============================================================================
// Purpose: Timer APB peripheral header
// Used in: cmsdk_apb_timer
//==============================================================================
// Timer reset macros
`define ARM_CTRL_RESET          4'h0
`define ARM_VALUE_RESET         32'h0000_0000
`define ARM_RELOAD_RESET        32'h0000_0000
`define ARM_INTCLEAR_RESET      1'b0